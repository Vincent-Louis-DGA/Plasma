---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_Program is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram_Program is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"000000400340ac033c0003243c0008000cac3c243c241400ac34243c243c273c",
INIT_01 => X"00008c8c8c3caf00af00af2340afafafafafafafafafafafafafafafafafaf23",
INIT_02 => X"acacacac40033423038f038f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f23",
INIT_03 => X"000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403acacacacacacacac",
INIT_04 => X"0000afafafaf272703008f240c3c000caf2700030014009024ac303c00100090",
INIT_05 => X"00a024008c001030008d343c353c001827038f8f8f8f02021402260c9002001a",
INIT_06 => X"8c343c301030008c343c30038c343c1030008c343c3c1430008c343c00030014",
INIT_07 => X"00030000109000900010001400240010001400900090000018ac033c00143000",
INIT_08 => X"1400240024241000102c0090000018000003a00024140090a000249000100090",
INIT_09 => X"0300140000240000002490000018000003001400002400249000001800000300",
INIT_0A => X"001000900010ad0014009024140090ad24248d00142c2424100090ad00af2700",
INIT_0B => X"2414009000102c14002c242c0090241000140024100014009024142400242424",
INIT_0C => X"00142c24002703008f240c240010000c0011000010240c24241524ad00008d24",
INIT_0D => X"a02524a024042414a02590000000000000000000143c142400001400243ca010",
INIT_0E => X"2400900030000000243c242424a024a02401030014002424a0a0909000100024",
INIT_0F => X"0caf27ac03af24343c8fac343ca003a09000309000243c00300003a000a00424",
INIT_10 => X"af272703008f00142824ac343c00240424ac2424acac00ac00ac00343c00af00",
INIT_11 => X"008c0010008ca00390ac008cac008c2703008f240c0010240c3c001428ac343c",
INIT_12 => X"27af0c24243c8e00afaf2700032400140090241000900014008c0010008c0014",
INIT_13 => X"2703008f240caf2727038f8f240caf278eaf14008f8e240c243c14343c8f240c",
INIT_14 => X"2703008f240caf272703008f240caf272703008f240caf272703008f240caf27",
INIT_15 => X"3002343c8c02343c1030008c022424243c363c00afafafafafafafafafafaf27",
INIT_16 => X"023c14003c8e3c102c1024001000100010001000920210270c02020c02001424",
INIT_17 => X"10020c0210020c0014000210020c0014000210020c001400920210270c02020c",
INIT_18 => X"afaf2727038f8f8f8f8f8f8f8f8f8fac008f8f02142e26ac02020c0202143402",
INIT_19 => X"2703008f8f8f008f020c02278f0000020c02278f0000020c27008f270c00afaf",
INIT_1A => X"2727038f8f8f8f260c0232a2260c3000a2260c3000a224000c0000afafafaf27",
INIT_1B => X"001030002703008fac0c248fac248fac243c8fac343cac343ca43ca43ca43caf",
INIT_1C => X"30ac3c3ca43ca43c24afaf27a4033ca43ca43c30030000003024140000302494",
INIT_1D => X"0c0032002400320000afafaf2727038f8fa6240c343cac3cac3ca6363ca43c34",
INIT_1E => X"3c8f8f8f300c26343c24140024a02430001826343ca43ca43c24a43ca43c2400",
INIT_1F => X"028fa6a626a6a6320c26000024323200000000363cafafafafaf8faf272703a4",
INIT_20 => X"ac3cac3cac3cac3cac3cac3cac343c343c000c003400afaf2727038f8f8f8f8f",
INIT_21 => X"a0240024a0240024a4240024ac00343c240424a0002424a43c24a43c24a43c24",
INIT_22 => X"3c363c3c00af343ca0acac243cafafafafafafaf2727038f8f240c242400af24",
INIT_23 => X"ae008f000caf2400008f001430008c343c1030008e240c26240c27270c8f2436",
INIT_24 => X"8f8f240c243c240c27270c001000102a260014282424142410002400343c00ae",
INIT_25 => X"8f00a0243c240c3c240c3424000c240c2424afafafafafafaf2727038f8f8f8f",
INIT_26 => X"0002af8f24140024a000343c24001430008c343c1030008eac24363c34363cac",
INIT_27 => X"343c0000000000000000000c000c270cafafaf27001000142eaeae00300c2602",
INIT_28 => X"0c26243c240cac24343cac243c343cac343c8c0000000000000000ae26363c8c",
INIT_29 => X"0c241400922410240c3c02020c00afafaf270010320c00000c270c240c2702ae",
INIT_2A => X"8c00343cafafafaf2727038f8f8f020c0010020c0014000010020c2414001002",
INIT_2B => X"003c8e3c102c1024001000102410241000922410240c3c02020c020014243000",
INIT_2C => X"0010020c0014000010020c24140010020c241400922410240c3c02020c023c14",
INIT_2D => X"31333742464a4e52565a0a00000000000027038f8f8f8f020c0014340010020c",
INIT_2E => X"01000000726f48363131310a70446f4421630a00433834305854504c48443935",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000020202020",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"00000084e00244e00200e042020000000062034202a560a4a01d8404a5059c1c",
INIT_01 => X"a086c6c5c406bb00bb00ba5a1abfb9b8afaeadacabaaa9a8a7a6a5a4a3a2a1bd",
INIT_02 => X"939291909b401bbd60bb60bbbabfb9b8afaeadacabaaa9a8a7a6a5a4a3a2a1a5",
INIT_03 => X"00e000c4e0000085a2e09f9d9c9e979695949392919002e09f9d9c9e97969594",
INIT_04 => X"a000b0b1b2bfbdbde000bf8400040000bfbd00e0004000828462420300400082",
INIT_05 => X"c543c686e30040420002e707080800a0bde0b0b1b2bf20504011100044508020",
INIT_06 => X"6263038440420042420242e042420240420062630302404200424202c0e00040",
INIT_07 => X"00e000620042a74387e68740e6e7006000620042a7438700c044e00200404200",
INIT_08 => X"40e5e743424200064062004387e0a000c0e04086c64000a26286a5a2004000a2",
INIT_09 => X"e00040e54342024606e74387e0a000e0e00040c5434207c64386c0a000c0e000",
INIT_0A => X"00400062000020854000824240008222428422004042420840008220a0bfbdc0",
INIT_0B => X"a54000e20040c2606242c2c300e60800004a000800004b0082e7aca5600a0b0c",
INIT_0C => X"004042c2a0bde000bfa50084000000000002000000a5008402020222450022a5",
INIT_0D => X"e008e7e20261e780e20842496b008600000006008101c1010786c0804902a000",
INIT_0E => X"e7a7636863c383c94802090607a202a20200e00040a7a5e7a3e2e3a20040a7e7",
INIT_0F => X"00bfbd62e08242630382444202a2e0a6828384464363030282e0e040a743c1c6",
INIT_10 => X"bfbdbde000bf0040a2a56563030042a1a5454205858305830583058404408200",
INIT_11 => X"0082006000a3a2e082a20082a20082bde000bf84000000840004004082444202",
INIT_12 => X"a4a2000584040280b0bfbd00e00200a3008302a000a500620082006000a30062",
INIT_13 => X"bde000bf0400bfbdbde0b0bf0500828402a24300830205008404436303a20500",
INIT_14 => X"bde000bf0400bfbdbde000bf0400bfbdbde000bf0400bfbdbde000bf0400bfbd",
INIT_15 => X"432363034222420240420042341516171e941400a4b0b1b2b3b4b5b6b7bebfbd",
INIT_16 => X"0002438203040240826202000000550056005700423440c50040400000606202",
INIT_17 => X"000000340000000055003400000000560034000000005700623440c500606000",
INIT_18 => X"b2bfbdbde0b0b1b2b3b4b5b6b7bebf4600a68234402231403420000034824234",
INIT_19 => X"bde062b0b1b212bf300002a5a26212300002a5a262123000a540b0a50080b0b1",
INIT_1A => X"bdbde0b0b1b2bf05002031120500841112050084111212a0001180b0b1b2bfbd",
INIT_1B => X"60a0a500bde000bf4000048262028362420283404202404202260125012401bf",
INIT_1C => X"a52201022401220102b0bfbd26e0012501240142e0066206c3844065c2636382",
INIT_1D => X"006010e005a024c080b0b1bfbdbde0b0bf0205008404270126010010102501a5",
INIT_1E => X"01b0b1bfa5002584048440656382426200a02584043001220102200122010240",
INIT_1F => X"80bf60725271708400546040053110e0c0a0807313b0b1b3b4bfb2b2bdbde022",
INIT_20 => X"200120012001200120013001a24202a5058000800480b0bfbdbde0b0b1b2b3b4",
INIT_21 => X"6202a4846202a4846202a48443a4630384616340a40304220102220102220102",
INIT_22 => X"1231111400824202604060430280b0b1b2b3b4bfbdbde0b0bf0700060500a484",
INIT_23 => X"4340840000824240008200404200626303404200220500840500a4a500841352",
INIT_24 => X"b4bf050084040500a4a5000080004002100040a2a563806340c36300c6060033",
INIT_25 => X"824080640384000406000504000006000504b0b1b2b3b4b5bfbdbde0b0b1b2b3",
INIT_26 => X"0060a58484406563830084040500404200626303404200228214521215311160",
INIT_27 => X"4202000000000000000000000000a400b0b1bfbd0000004002344540e7001015",
INIT_28 => X"0031840404006202630362420263034042025100000000000000001131101051",
INIT_29 => X"00028200240240a5000520200080b0b1bfbd00002400400000a4000600a52011",
INIT_2A => X"42a24202b0b1b2bfbdbde0b0b1bf000000000000008200000000000282000000",
INIT_2B => X"8203040240826202000000820282028200240240a50005202000006062024380",
INIT_2C => X"0000000000820000000000028200000000028200440240a50005404000000243",
INIT_2D => X"3232364145494d5155590d000000000000bde0b0b1b2bf000000824200000000",
INIT_2E => X"000000006c206534303639000a480a480a6b5300443935315955514d49454136",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"00000060006000002000001700000000040020000000ff180080170017009700",
INIT_01 => X"f8200000002000d800d800ff70000000000000000000000000000000000000ff",
INIT_02 => X"0000000060000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000201000000000000000000000000000000000000000000000000000",
INIT_04 => X"888000000000ff00000000160000000000ff000000ff00000000002000000000",
INIT_05 => X"100000100000000000000020002030000000000000001010ff10000000109000",
INIT_06 => X"000020000000000000200000000020ff000000002020000000000020100000ff",
INIT_07 => X"0000101000001000100010ff1000000000000000100010380000002000ff0000",
INIT_08 => X"ff100030ffff001100000000103000381000001000ff00000018000030000000",
INIT_09 => X"0000ff1030ff101010000010300038100000ff1038ff10000010380030100000",
INIT_0A => X"0000000010000018000000ffff000000000000000000ff00002800004800ff10",
INIT_0B => X"00ff0000000000001800ff000000000000000000000000000000000038000000",
INIT_0C => X"400000ff3800000000ff0100000000010000000000ff010000000000100000ff",
INIT_0D => X"00000000000000ff000000101058000000200000008000ff0000001816000000",
INIT_0E => X"0010001800181818170000000000000000100000ff1000ff00000000000010ff",
INIT_0F => X"0000ff000080000020800000200000000020000010170011001000001000ffff",
INIT_10 => X"00ff0000000000ff000000002028ffffff00010000001a001c001e0020288000",
INIT_11 => X"0000000000000000000000000000000000000000020000170000000000000020",
INIT_12 => X"00000000170000800000ff000000100000000000000010000000000000001000",
INIT_13 => X"00000000000000ff000000000000808000000000800000001700000000000000",
INIT_14 => X"00000000000000ff00000000000000ff00000000000000ff00000000000000ff",
INIT_15 => X"ff8040200010502000ff000010000000005020880000000000000000000000ff",
INIT_16 => X"200000104000f000060008000000000000000000001000170220280220200008",
INIT_17 => X"0020021000200200000010002002000000100020020000000010001702202802",
INIT_18 => X"0000ff0000000000000000000000000000008010ff0808001028022010000810",
INIT_19 => X"0000100000001a002001800000901a2001800000901a20010090000001880000",
INIT_1A => X"ff000000000000000120000000010022000001002400008001268800000000ff",
INIT_1B => X"3000ff180000000000000080000080000a008000582000502000200020002000",
INIT_1C => X"8020206d20202020450000ff30002030203020ff00103014ff00ff1030ff0000",
INIT_1D => X"0330ff800010ff8818000000ff00000000000003202020202020002020202080",
INIT_1E => X"20000000ff03ff202000ff10000000001800ff20202020202000202020200838",
INIT_1F => X"10000000000000ff0300383000ffff88801810202000000000000000ff000020",
INIT_20 => X"2020202020202020202020200006012020300328ff800000ff00000000000000",
INIT_21 => X"0000180000001800003518000010536300ffff00100000202054202035202002",
INIT_22 => X"2030200080805435001700170080000000000000ff00000000000300ff200000",
INIT_23 => X"0018800004800020008000ff0000003020000000000000170000000003800030",
INIT_24 => X"000000001700000000000300ff0000000000ff0000ff0000ff10001886002800",
INIT_25 => X"80980017001703007203957080045403350200000000000000ff000000000000",
INIT_26 => X"3028008000ff1000001820200000ff00000030200000000000003020ea302017",
INIT_27 => X"00200000000000000000200200010004000000ff00ff00ff00000028ff030038",
INIT_28 => X"0000170000000000002000070000200000200000000000000000000000002000",
INIT_29 => X"0200000000000017020020280280000000ff00ff000088000000000001002000",
INIT_2A => X"0010502000000000ff0000000000200200002002000000000020020000000020",
INIT_2B => X"104000f00006000800000000000000000000000017020020280220200008ff80",
INIT_2C => X"0000200200000000002002000000002002000000000000170200202802200000",
INIT_2D => X"3331353944484c50545800000000000000000000000000200200000800002002",
INIT_2E => X"0000000064576c00343832000043004300657400454136325a56524e4a464237",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"0000000008004408000008a800001100ec4c005c0004fd2a0000a800a0007001",
INIT_01 => X"0924504c400060125c1058fc0054504c4844403c3834302c2824201c18141098",
INIT_02 => X"0c080400000801681360115c5854504c4844403c3834302c2824201c18141000",
INIT_03 => X"00080c000810121900082c2824201c1814100c08040000082c2824201c181410",
INIT_04 => X"25251014181ce018080010d48000008010e8000800fa00000100ff0000090000",
INIT_05 => X"2a00012100000808000004000800251120081014181c2521fb2a01d600212508",
INIT_06 => X"000800ff080100000800ff08000400fc080000080000080800000800250800f5",
INIT_07 => X"0008252302002100210621f52a01000500070000210021250e00080000fc0100",
INIT_08 => X"f32a0121c9d00200033a000021250f252508002101f900000021010025090000",
INIT_09 => X"0800f62a21d0402180010021250c25250800f82a21d040010021250a25250800",
INIT_0A => X"00220000253c0021040000d0f600000001010000090ad064122500002510e825",
INIT_0B => X"01e60000000647082507c6300000620b000300781000030001010c0125627801",
INIT_0C => X"250323fe2518080010fe230200040031000500000bfe100262067800210000ff",
INIT_0D => X"000101002d0401eb000123212312180000120d00020004ff0d1a0225d800002c",
INIT_0E => X"01210021ff06240420000f1c0201780030250800f82b01ff00000000000a2bff",
INIT_0F => X"1310e80008200160002000440001080000210f0021200002ff2508002100f6fc",
INIT_10 => X"10e81808001000fc640100600025fcfdff008c63000003000300036000253000",
INIT_11 => X"00000005000008080900000c04001018080010011e0003348000000665006000",
INIT_12 => X"1010990640001425181ce00008012502000801060008250a0004000500042512",
INIT_13 => X"1808001043d610e82008181c049928282c1006003420069948000e4344100499",
INIT_14 => X"1808001041d610e81808001049d610e81808001055d610e81808001054d610e8",
INIT_15 => X"ff260001002630014fff00002606011100200125381014181c2024282c3034c8",
INIT_16 => X"250123240000002e002d06002900270022001d0008263e743a25253125251300",
INIT_17 => X"082590260c258000050026132578000500261a2588000500082622743a252531",
INIT_18 => X"2024d838081014181c2024282c30340000381426a80100002625982526050026",
INIT_19 => X"280821181c20002421412110102100214121101021002141102510104125181c",
INIT_1A => X"e820081014181c09e725ff0806e7ff020503e7ff02022e25e702251014181ce0",
INIT_1B => X"2508ff2518080010001a011000041c008000180020010020012c012801240110",
INIT_1C => X"ff0401f302010001001014e82c080128012401ff08272102ff02fa2b21ff0200",
INIT_1D => X"9425ff250125ff2525101418e01808101400147c000110010c01000a01080100",
INIT_1E => X"01101418ff7cec140101fa2a0100610f2508e41c011a01180101160114010025",
INIT_1F => X"25240604080200ff941c252511ffff25252525140110141c20243818d8200816",
INIT_20 => X"340130012c012801240120010000011c01258d25ff25181ce028081014181c20",
INIT_21 => X"00ff210100012102000121040021638201fcff0021c9223c01413a014438010a",
INIT_22 => X"01000100253441440874047400282024282c3034c82008181c43e344ff251001",
INIT_23 => X"0025280007340125003400fc0400000001070400000199500b99101040280220",
INIT_24 => X"3034019950000b9910104000ce00030a0100f66401ff0501fe2a01259f012500",
INIT_25 => X"2825087400541d001f8d00f3254b415f440a181c2024282c30c838082024282c",
INIT_26 => X"2525102801fc2a0100251c011000fc0400000001070400000402200160000174",
INIT_27 => X"70000000000000000000251e00fd10a6505458a000ff00df20000025ffe30121",
INIT_28 => X"80016400011a00ff500000cc004c000040000000000000000000000001600000",
INIT_29 => X"88010500081118743a0025253125101418e000faffd62500c4108e0a9b102500",
INIT_2A => X"002630011014181ce02008101418259000032580000500000a25780605001025",
INIT_2B => X"240000002d002d06002900270622011e0008113c743a0025253125251400ff25",
INIT_2C => X"000a25800005000011257806050017258801050008111f743a00252531250123",
INIT_2D => X"3430343843474b4f53570000000000000020081014181c259800030000062590",
INIT_2E => X"00010100206f6c002e2e2e000050005000646100464237330057534f4b474338",
INIT_2F => X"00000000000000000000000000000000000000000000000000000000504c4440",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
