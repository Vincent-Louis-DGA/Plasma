---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_Program is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram_Program is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"00000040000340ac033c0003243c08000cac3c243c241400ac34243c243c273c",
INIT_01 => X"00008c8c8c3caf00af00af2340afafafafafafafafafafafafafafafafafaf23",
INIT_02 => X"acacacac40033423038f038f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f23",
INIT_03 => X"000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403acacacacacacacac",
INIT_04 => X"0000afafafaf272703008f240c3c000caf2700030014009024ac303c00100090",
INIT_05 => X"00a024008c001030008d343c353c001827038f8f8f8f02021402260c9002001a",
INIT_06 => X"8c343c301030008c343c30038c343c1030008c343c3c1430008c343c00030014",
INIT_07 => X"00030000109000900010001400240010001400900090000018ac033c00143000",
INIT_08 => X"1400240024241000102c0090000018000003a00024140090a000249000100090",
INIT_09 => X"0300140000240000002490000018000003001400002400249000001800000300",
INIT_0A => X"001000900010ad0014009024140090ad24248d00142c2424100090ad00af2700",
INIT_0B => X"2414009000102c14002c242c0090241000140024100014009024142400242424",
INIT_0C => X"00142c24002703008f240c240010000c0011000010240c24241524ad00008d24",
INIT_0D => X"a02524a024042414a02590000000000000000000143c142400001400243ca010",
INIT_0E => X"2400900030000000243c242424a024a02401030014002424a0a0909000100024",
INIT_0F => X"acac00ac00ac00343c00af000caf27ac03af24343c8fac343c0003a000a00424",
INIT_10 => X"0c0010240c3c001428ac343caf272703008f00142824ac343c00240424ac2424",
INIT_11 => X"001430008e00363c363c363c00a2a2a22400afafafafafafafaf272703008f24",
INIT_12 => X"0c020c262426a002240c02028e001030008c343c1430008eae001030008c343c",
INIT_13 => X"00000000000024028c343c020c240c3c000c00000000000024028c343c142a02",
INIT_14 => X"30008c343c1030008e363c363c363c1430008c343cac24343c020c240c3c000c",
INIT_15 => X"0000000c000c270cafafaf2727038f8f8f8f8f8f8f8f001030008e320c8e0014",
INIT_16 => X"343cac243c343cac343c8c0000000000000000ae26363c8c343c000000000000",
INIT_17 => X"52565a0a0000000000000010320c00000c270c240c2702ae0c26243c240cac24",
INIT_18 => X"0000726f486452645421630a00433834305854504c4844393531333742464a4e",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"0000008400e00244e00200e0420200000062034202a560a4a01d8404a5059c1c",
INIT_01 => X"a086c6c5c406bb00bb00ba5a1abfb9b8afaeadacabaaa9a8a7a6a5a4a3a2a1bd",
INIT_02 => X"939291909b401bbd60bb60bbbabfb9b8afaeadacabaaa9a8a7a6a5a4a3a2a1a5",
INIT_03 => X"00e000c4e0000085a2e09f9d9c9e979695949392919002e09f9d9c9e97969594",
INIT_04 => X"a000b0b1b2bfbdbde000bf8400040000bfbd00e0004000828462420300400082",
INIT_05 => X"c543c686e30040420002e707080800a0bde0b0b1b2bf20504011100044508020",
INIT_06 => X"6263038440420042420242e042420240420062630302404200424202c0e00040",
INIT_07 => X"00e000620042a74387e68740e6e7006000620042a7438700c044e00200404200",
INIT_08 => X"40e5e743424200064062004387e0a000c0e04086c64000a26286a5a2004000a2",
INIT_09 => X"e00040e54342024606e74387e0a000e0e00040c5434207c64386c0a000c0e000",
INIT_0A => X"00400062000020854000824240008222428422004042420840008220a0bfbdc0",
INIT_0B => X"a54000e20040c2606242c2c300e60800004a000800004b0082e7aca5600a0b0c",
INIT_0C => X"004042c2a0bde000bfa50084000000000002000000a5008402020222450022a5",
INIT_0D => X"e008e7e20261e780e20842496b008600000006008101c1010786c0804902a000",
INIT_0E => X"e7a7636863c383c94802090607a202a20200e00040a7a5e7a3e2e3a20040a7e7",
INIT_0F => X"85830583058305840440820000bfbd62e08242630382444202e0e040a743c1c6",
INIT_10 => X"000000840004004082444202bfbdbde000bf0040a2a56563030042a1a5454205",
INIT_11 => X"1140420062409414b5157313004242420280b0b1b2b3b4b5b6bfbdbde000bf84",
INIT_12 => X"000000310645564206004020900040420062630340420062a211404200626303",
INIT_13 => X"9004900490100640504202400084000404009004900490100640504202402240",
INIT_14 => X"4200626303404200623111521273134042004242026202630340008400040400",
INIT_15 => X"000000000000a400b0b1bfbdbde0b0b1b2b3b4b5b6bf00404200220400500040",
INIT_16 => X"6303624202630340420251000000000000000011311010514202000000000000",
INIT_17 => X"5155590d00000000000000002400400000a4000600a520110031840404006202",
INIT_18 => X"00006c2065207820780a6b5300443935315955514d494541363232364145494d",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"0000006000006000002000000c000000020020000000ff1800800c000c008c00",
INIT_01 => X"f8200000002000d800d800ff70000000000000000000000000000000000000ff",
INIT_02 => X"0000000060000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000201000000000000000000000000000000000000000000000000000",
INIT_04 => X"888000000000ff000000000b0000000000ff000000ff00000000002000000000",
INIT_05 => X"100000100000000000000020002030000000000000001010ff10000000109000",
INIT_06 => X"000020000000000000200000000020ff000000002020000000000020100000ff",
INIT_07 => X"0000101000001000100010ff1000000000000000100010380000002000ff0000",
INIT_08 => X"ff100030ffff001100000000103000381000001000ff00000018000030000000",
INIT_09 => X"0000ff1030ff101010000010300038100000ff1038ff10000010380030100000",
INIT_0A => X"0000000010000018000000ffff000000000000000000ff00002800004800ff10",
INIT_0B => X"00ff0000000000001800ff000000000000000000000000000000000038000000",
INIT_0C => X"400000ff3800000000ff0100000000010000000000ff010000000000100000ff",
INIT_0D => X"00000000000000ff000000101058000000200000008000ff000000180b000000",
INIT_0E => X"00100018001818180c0000000000000000100000ff1000ff00000000000010ff",
INIT_0F => X"00001a001c001e00202880000000ff000080000020800000201000001000ffff",
INIT_10 => X"0200000c000000000000002000ff0000000000ff000000002028ffffff000100",
INIT_11 => X"1600000000b00020002000208800000000900000000000000000ff0000000000",
INIT_12 => X"0020010000000010000128200000ff0000000020000000000016ff0000000020",
INIT_13 => X"202120202020002800002020000c000021012021202020200028000020ff0020",
INIT_14 => X"0000000020000000000020002000200000000000200000002020000c00002101",
INIT_15 => X"0000200200010002000000ff0000000000000000000000ff00000000000000ff",
INIT_16 => X"0020000700002000002000000000000000000000000020000020000000000000",
INIT_17 => X"5054580000000000000000ff00008800000000000100200000000c0000000000",
INIT_18 => X"000064576c0050005000657400454136325a56524e4a4642373331353944484c",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"00000000000800440800000884001100b44c00580004fd2a0000840080006901",
INIT_01 => X"0924504c400060125c1058fc0054504c4844403c3834302c2824201c18141098",
INIT_02 => X"0c080400000801681360115c5854504c4844403c3834302c2824201c18141000",
INIT_03 => X"00080c000810121900082c2824201c1814100c08040000082c2824201c181410",
INIT_04 => X"25251014181ce018080010f08000008010e8000800fa00000100ff0000090000",
INIT_05 => X"2a00012100000808000004000800251120081014181c2521fb2a01d600212508",
INIT_06 => X"000800ff080100000800ff08000400fc080000080000080800000800250800f5",
INIT_07 => X"0008252302002100210621f52a01000500070000210021250e00080000fc0100",
INIT_08 => X"f32a0121c9d00200033a000021250f252508002101f900000021010025090000",
INIT_09 => X"0800f62a21d0402180010021250c25250800f82a21d040010021250a25250800",
INIT_0A => X"00220000253c0021040000d0f600000001010000090ad064122500002510e825",
INIT_0B => X"01e60000000647082507c6300000620b000300781000030001010c0125627801",
INIT_0C => X"250323fe2518080010fe230200040031000500000bfe100262067800210000ff",
INIT_0D => X"000101002d0401eb000123212312180000120d00020004ff0d1a0225f400002c",
INIT_0E => X"01210021ff0624043c000f1c0201780030250800f82b01ff00000000000a2bff",
INIT_0F => X"0000030003000360002517001210e8000813016000130044002508002100f6fc",
INIT_10 => X"12000350800000066500600010e81808001000fc640100600025fcfdff008c63",
INIT_11 => X"000801000025080104010c012502010020251014181c2024282cd01808001001",
INIT_12 => X"8e259b0110030021109b25250000fc0100000c01070100000000fc0100000c01",
INIT_13 => X"210023c021800a25001401258e5c8000439b210023c021800a25001001d80225",
INIT_14 => X"0200000c0107020000080020010c0119010000080000080c01258e648000439b",
INIT_15 => X"0000251200f11025505458a030081014181c2024282c00ee010000ffd60000fc",
INIT_16 => X"5000009c004c0000400000000000000000000000016000007000000000000000",
INIT_17 => X"4f53570000000000000000faffd62500c4108e0a9b10250080016c00011900ff",
INIT_18 => X"0000206f6c0072007200646100464237330057534f4b4743383430343843474b",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
