---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_PlasmaBootLoader is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram_PlasmaBootLoader is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"afafafafafafafafaf23ac033c08000cac3c243c241400ac273c243c243c273c",
INIT_01 => X"8f8f8f8f8f8f8f8f8f2300008c8c8c3caf00af00af2340afafafafafafafafaf",
INIT_02 => X"acacacacacacacacacacac40034040033423038f038f8f8f8f8f8f8f8f8f8f8f",
INIT_03 => X"ac303c00100090000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403ac",
INIT_04 => X"02260c9002001a0000afafafaf272703008f240c3c000caf2700030014009024",
INIT_05 => X"8c343c0003001400a024008c001030008d343c353c001827038f8f8f8f020214",
INIT_06 => X"ac033c001430008c343c301030008c343c30038c343c1030008c343c3c143000",
INIT_07 => X"0024900010009000030000109000900010001400240010001400900090000018",
INIT_08 => X"000018000003001400240024241000102c0090000018000003a00024140090a0",
INIT_09 => X"0090ad00af270003001400002400000024900000180000030014000024002490",
INIT_0A => X"24142400242424001000900010ad0014009024140090ad24248d00142c242410",
INIT_0B => X"1524ad00008d242414009000102c14002c242c00902410001400241000140090",
INIT_0C => X"001400243ca01000142c24002703008f240c240010000c0011000010240c2424",
INIT_0D => X"a0909000100024a02524a024042414a02590000000000000000000143c142400",
INIT_0E => X"0003a000a004242400900030000000243c242424a024a02401030014002424a0",
INIT_0F => X"243c353c00243c18ac000001343c01009000243cac03343c24042424ac24343c",
INIT_10 => X"140024ad242404240030002490adad0000912590001400009100243c24353c00",
INIT_11 => X"1800002703008f240c2700a3a300a300af272703008f240c2700a3af27000300",
INIT_12 => X"14002400a0000014303000300000ac8d240424acad2424353c24343c24353c00",
INIT_13 => X"020c02020c323200000000afafafafafaf8faf8faf8faf27ac0324343c000324",
INIT_14 => X"afafaf8f2727038f8f8f8f8f8f8f8f8f000c020c8f021a020c02021a020c021a",
INIT_15 => X"8f000c00240000afaf272703008faf0cafafafaf308f272703008faf0c0030af",
INIT_16 => X"af24afaf272703008f000c000024afaf272703008f000c000024afaf27270300",
INIT_17 => X"000024af24af2727030000000000008f8f93939393270c000024af270c000024",
INIT_18 => X"1a240c3c270c240c2702000c00243c00afafafafafaf27270300008f9393270c",
INIT_19 => X"8f8f8f8f8f240c3c02140226260c001032270c260c001028240c2790023c3c00",
INIT_1A => X"3cafaf2727038f8f240c2702270c000224af24240424a0272400afaf2727038f",
INIT_1B => X"0c2792240c8e000c92263cafaf2727038f8f93000c240c2792240c8e000c9226",
INIT_1C => X"af2727038f8f93000c240c2792240c8e000c92263cafaf2727038f8f93000c24",
INIT_1D => X"14002c2c3830a3af0cafaf272703008f000c0010243000000c0010243000000c",
INIT_1E => X"00000024afafaf2493af0c008c0000263c000024afafaf93a324a32424142424",
INIT_1F => X"af2727038f8f8fa30010a32414240010a32410002c2c3830a3000caf0c278c00",
INIT_20 => X"0c270c02000c243c000c270c270c02000c243c000c270c270c02000c243caf0c",
INIT_21 => X"0c3cafaf2727038f8f270c270c02240c3c00000c270c270c02240c3c00000c27",
INIT_22 => X"000c000c000caf272703248f8f240c273c270c000024af24020c240c02279324",
INIT_23 => X"0c273c000caf27ac03343cac24343cac343c2703008f3c0c340c3c340c3c3c0c",
INIT_24 => X"02142a26ae0000000c3c0200afafafaf272703008f240c003caf3c240c273c24",
INIT_25 => X"000c363c001aaeafae0c00ae0c24363cac24343cafafafafaf2727038f8f8f8f",
INIT_26 => X"8e363cac24343cafafaf2727038f8f8f8f8fac0c24343c00140226ac00008fae",
INIT_27 => X"565a0a0000000000002703008f8fac0024343c10008f000c0010000c00103000",
INIT_28 => X"523220523100203020205200433834305854504c4844393531333742464a4e52",
INIT_29 => X"00000000000000000000ff0807070e01000000000000734c204e205620523420",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"a9a8a7a6a5a4a3a2a1bd44e00200000062034202a560a4a0bd1d8404a5059c1c",
INIT_01 => X"a9a8a7a6a5a4a3a2a1a5a086c6c5c406bb00bb00ba5a1abfb9b8afaeadacabaa",
INIT_02 => X"9d9c9e979695949392919084e0029b401bbd60bb60bbbabfb9b8afaeadacabaa",
INIT_03 => X"6242030040008200e000c4e0000085a2e09f9d9c9e979695949392919002e09f",
INIT_04 => X"11100044508020a000b0b1b2bfbdbde000bf8400040000bfbd00e00040008284",
INIT_05 => X"424202c0e00040c543c686e30040420002e707080800a0bde0b0b1b2bf205040",
INIT_06 => X"44e002004042006263038440420042420242e042420240420062630302404200",
INIT_07 => X"86a5a2004000a200e000620042a74387e68740e6e7006000620042a7438700c0",
INIT_08 => X"86c0a000c0e00040e5e743424200064062004387e0a000c0e04086c64000a262",
INIT_09 => X"008220a0bfbdc0e00040e54342024606e74387e0a000e0e00040c5434207c643",
INIT_0A => X"e7aca5600a0b0c00400062000020854000824240008222428422004042420840",
INIT_0B => X"020222450022a5a54000e20040c2606242c2c300e60800004a000800004b0082",
INIT_0C => X"86c0804902a000004042c2a0bde000bfa50084000000000002000000a5008402",
INIT_0D => X"e2e3a20040a7e7e008e7e20261e780e20842496b008600000006008101c10107",
INIT_0E => X"e0e040a743c1c6e7a7636863c383c94802090607a202a20200e00040a7a5e7a3",
INIT_0F => X"42028c0cc24202a062c505406303400042c2420240e042024241420262026303",
INIT_10 => X"40e5e7206363616340424803c22e824800624a488a40e200a2c242020e2909c2",
INIT_11 => X"a00500bde000bf0500a4a0a4a204a204bfbdbde000bf0500a4a0a4bfbd00e000",
INIT_12 => X"40c5c6004382064ac24343420203e002424142eb2c020a08080be7070c290960",
INIT_13 => X"40000060005310e0c0a080b0b1b3b4b5bfb7b7b6b6b2b2bd62e002630300e002",
INIT_14 => X"a7a0bfa2bdbde0b0b1b2b3b4b5b6b7bf00006000a4e0e04000c0a0c040008020",
INIT_15 => X"bf80004004a080a6bfbdbde000bfa200a0a0a0bf84a2bdbde000bfa2000084a0",
INIT_16 => X"b010b0bfbdbde000bfa000a00004a0bfbdbde000bfa000a00004a0bfbdbde000",
INIT_17 => X"a00004a202bfbdbde0454404430302b0bfa5a4a3a2a700a00004b0a700a00004",
INIT_18 => X"20840004a4000600a500c000a0840480b0b1b2b3b4bfbdbde04302bfa3a2a700",
INIT_19 => X"b1b2b3b4bf840004904011104400004002a40064000040420600a54490121300",
INIT_1A => X"10b0bfbdbde0b0bf0600a500a700800004a20242616340a20380b0bfbdbde0b0",
INIT_1B => X"00a4060400050000041010b0bfbdbde0b0bfa200000500a40604000500000410",
INIT_1C => X"bfbdbde0b0bfa200000500a4060400050000041010b0bfbdbde0b0bfa2000005",
INIT_1D => X"40438342824482b000b1bfbdbde000bf00008062024340000080620283400000",
INIT_1E => X"02a00004a0a0b11182a200a04250021010a00004a0a0a082a202820202820202",
INIT_1F => X"bfbdbde0b0b1bf9100008202820200008202404383428244820000a200a74250",
INIT_20 => X"00a50000400084040000a400a50000400084040000a400a5000040008404b000",
INIT_21 => X"0004b0bfbdbde0b0bfa400a50000840004400000a400a50000840004400000a4",
INIT_22 => X"000000000000bfbdbde002b0bf0600a504a700a00004a2020000060000b08484",
INIT_23 => X"00a5040000bfbd44e0420262026303404202bde000bf04008400048400040400",
INIT_24 => X"004022315062100000120000b0b1b2bfbdbde000bf0600400482020600a50406",
INIT_25 => X"0000731300400282120040020002101062026303b0b1b2b3bfbdbde0b0b1b2bf",
INIT_26 => X"0210106202630380b0bfbdbde0b0b1b2b3bf6200026303004032317071408371",
INIT_27 => X"55590d000000000000bde000b0bf628002630380008400000000000000404200",
INIT_28 => X"20560020560000003a006500443935315955514d494541363232364145494d51",
INIT_29 => X"00000000000000000000ff0406030c0200000000000020693a563a4300205600",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000ff0000200000040020000000ff18001600160014009400",
INIT_01 => X"00000000000000000000f8200000002000d800d800ff70000000000000000000",
INIT_02 => X"0000000000000000000000600060600000000000000000000000000000000000",
INIT_03 => X"0000200000000000000000002010000000000000000000000000000000000000",
INIT_04 => X"10000000109000888000000000ff00000000130000000000ff000000ff000000",
INIT_05 => X"000020100000ff100000100000000000000020002030000000000000001010ff",
INIT_06 => X"00002000ff0000000020000000000000200000000020ff000000002020000000",
INIT_07 => X"180000300000000000101000001000100010ff10000000000000001000103800",
INIT_08 => X"10380030100000ff100030ffff001100000000103000381000001000ff000000",
INIT_09 => X"2800004800ff100000ff1030ff101010000010300038100000ff1038ff100000",
INIT_0A => X"000000380000000000000010000018000000ffff000000000000000000ff0000",
INIT_0B => X"000000100000ff00ff0000000000001800ff0000000000000000000000000000",
INIT_0C => X"00001813000000400000ff3800000000ff0100000000010000000000ff010000",
INIT_0D => X"000000000010ff00000000000000ff000000101058000000200000008000ff00",
INIT_0E => X"1000001000ffff0010001800181818140000000000000000100000ff1000ff00",
INIT_0F => X"140000206814000000282838002040500010140000000020ffffff0000000020",
INIT_10 => X"ff10000000ffffff400010000000001000000000100010000030140000002058",
INIT_11 => X"0028180000000000010030000012001400ff00000000000100300000ff000000",
INIT_12 => X"ff100018001010000000100010180000ffffff00000000002000002000002030",
INIT_13 => X"28022020010000a888a080000000000000000000000000ff0000000020000000",
INIT_14 => X"00000000ff000000000000000000000000023002002800300128200028022000",
INIT_15 => X"003002280038100000ff000000000002000000000000ff000000000002380000",
INIT_16 => X"00000000ff0000000038023028000000ff0000000038023028000000ff000000",
INIT_17 => X"302800000000ff0000101022101c160000000000000002302800000002302800",
INIT_18 => X"001400000000000100208800a0140080000000000000ff000010120000000002",
INIT_19 => X"000000000014000010ff10001400000000000014000000000001000010000080",
INIT_1A => X"000000ff000000000003002000023028000000ffffff000000800000ff000000",
INIT_1B => X"02000000020000010014000000ff000000000000020002000000020000010014",
INIT_1C => X"00ff000000000000020002000000020000010014000000ff0000000000000200",
INIT_1D => X"0010000000008000030000ff0000000000031000000020000310000000200003",
INIT_1E => X"1030280000000000800002380010101400302800000000800000800000000000",
INIT_1F => X"00ff000000000080000080000000000080000010000000008000030002000010",
INIT_20 => X"0000012080001400000300000001208000140000030000000120800014000003",
INIT_21 => X"00000000ff000000000000000120140000800002000000012014000080000200",
INIT_22 => X"00030004000300ff00000000000003001d000230280000002000000128008014",
INIT_23 => X"020000000300ff00000020000000200000200000000000030103000003000003",
INIT_24 => X"10ff000000801a000020888000000000ff000000000702280080400003000000",
INIT_25 => X"00040020880000800004900004000020000000200000000000ff000000000000",
INIT_26 => X"00002000000020800000ff00000000000000000000002000ff10000018808000",
INIT_27 => X"545800000000000000000010000000f8000020ff008000040000000400000000",
INIT_28 => X"204500204500000020006100454136325a56524e4a4642373331353944484c50",
INIT_29 => X"000000000000000000000102040100040000000000003a6e2043205200204500",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"302c2824201c181410984408001200d54c004c0004fd2a00c800e000d800c301",
INIT_01 => X"302c2824201c181410000924504c400060125c1058fc0054504c4844403c3834",
INIT_02 => X"2824201c1814100c080400000800000801681360115c5854504c4844403c3834",
INIT_03 => X"00ff000009000000080c000810121900082c2824201c1814100c08040000082c",
INIT_04 => X"2a01cf0021250825251014181ce018080010f47900007910e8000800fa000001",
INIT_05 => X"000800250800f52a00012100000808000004000800251120081014181c2521fb",
INIT_06 => X"00080000fc0100000800ff080100000800ff08000400fc080000080000080800",
INIT_07 => X"210100250900000008252302002100210621f52a01000500070000210021250e",
INIT_08 => X"21250a25250800f32a0121c9d00200033a000021250f252508002101f9000000",
INIT_09 => X"2500002510e8250800f62a21d0402180010021250c25250800f82a21d0400100",
INIT_0A => X"010c012562780100220000253c0021040000d0f600000001010000090ad06412",
INIT_0B => X"067800210000ff01e60000000647082507c6300000620b000300781000030001",
INIT_0C => X"1a0225f800002c250323fe2518080010fe1c020004002a000500000bfe090262",
INIT_0D => X"000000000a2bff000101002d0401eb000123212312180000120d00020004ff0d",
INIT_0E => X"2508002100f6fc01210021ff06240440000f1c0201780030250800f82b01ff00",
INIT_0F => X"cc00c40021c800280007c025c80025250021c4000008c000ffffff010002c000",
INIT_10 => X"e72a010001ffffff25ff04010000000700000100210324000021c00001c00021",
INIT_11 => X"21c0252008001803ec1025121103100318e02008001801ec10251018e0000800",
INIT_12 => X"eb2a01250021c30407ff210142400000ffffff00000107c40001c0000fc80025",
INIT_13 => X"25232525e0ffff2525252510141c202430502c48285418c8000802c000000801",
INIT_14 => X"14102038d838081014181c2024282c300063253d4c250425ec252504252e2503",
INIT_15 => X"18259b250325251018e02808002010681c181420ff38d828080020186825ff1c",
INIT_16 => X"10022024d82008001825a92525041018e02008001825a92525061018e0200800",
INIT_17 => X"2525b5100220d8280825210021000020241b1a19181a9b25256510189b252585",
INIT_18 => X"185c79001079109410252579255400255054585c60649828082500201918189b",
INIT_19 => X"54585c606468870021ed2a016479000301107960790003021094100021000025",
INIT_1A => X"00181ce03808303414091825189b2525031014fffdff002b13253034c8680850",
INIT_1B => X"3d100b65230800e00bac00181ce02008181c100063013d100765230400e007ac",
INIT_1C => X"10e82008181c100063013d101365231000e013ac00181ce02008181c10006301",
INIT_1D => X"0525010140e011289e2c30c818080010005c250380c0250072250ac0c025005c",
INIT_1E => X"8025256118141001131c6825002180ac002525061814101320ff130201028004",
INIT_1F => X"54a83808282c3013000213020480000813040425010140e011009e1c68200021",
INIT_20 => X"8710c825257984000088108710c825257978000072108710c82525796c00505c",
INIT_21 => X"790070748858085054108710c8259879002500f9108710c8259079002500db10",
INIT_22 => X"00fe003b00b410e8780801707414091800189b25259f101425870a94253013a0",
INIT_23 => X"b6102000b418e00008400000fa80000094001808001020430043181043181843",
INIT_24 => X"25f8040100210000bd0025251014181ce02008001800b6252019000809102008",
INIT_25 => X"008f6000250e0019008f25008f2a6000000110001014181c20d820081014181c",
INIT_26 => X"00740000546000191014e828081014181c2000bdff600000f62a040021251900",
INIT_27 => X"53570000000000000018082510140009ff6000f200190079000300a600050800",
INIT_28 => X"3a43003a4300000000006400464237330057534f4b4743383430343843474b4f",
INIT_29 => X"00000000000000000000000000000000020001000000206500520020003a4300",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
