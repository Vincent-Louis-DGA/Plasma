---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_Program is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram_Program is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"afafafafafafafafaf23ac033c08000cac3c243c241400ac273c243c243c273c",
INIT_01 => X"8f8f8f8f8f8f8f8f8f2300008c8c8c3caf00af00af2340afafafafafafafafaf",
INIT_02 => X"acacacacacacacacacacac40034040033423038f038f8f8f8f8f8f8f8f8f8f8f",
INIT_03 => X"ac303c00100090000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403ac",
INIT_04 => X"02260c9002001a0000afafafaf272703008f240c3c000caf2700030014009024",
INIT_05 => X"8c343c0003001400a024008c001030008d343c353c001827038f8f8f8f020214",
INIT_06 => X"ac033c001430008c343c301030008c343c30038c343c1030008c343c3c143000",
INIT_07 => X"0024900010009000030000109000900010001400240010001400900090000018",
INIT_08 => X"000018000003001400240024241000102c0090000018000003a00024140090a0",
INIT_09 => X"0090ad00af270003001400002400000024900000180000030014000024002490",
INIT_0A => X"24142400242424001000900010ad0014009024140090ad24248d00142c242410",
INIT_0B => X"1524ad00008d242414009000102c14002c242c00902410001400241000140090",
INIT_0C => X"001400243ca01000142c24002703008f240c240010000c0011000010240c2424",
INIT_0D => X"a0909000100024a02524a024042414a02590000000000000000000143c142400",
INIT_0E => X"0003a000a004242400900030000000243c242424a024a02401030014002424a0",
INIT_0F => X"3c24363c373c363c24ac343c00afafafafafafafafafaf270003001c00300018",
INIT_10 => X"008f001430008e00100000001200aeac3caf0c343c8c343cae24360236023c36",
INIT_11 => X"001430008e001430008c24a000008f0010288e343c001030008eaeae24009000",
INIT_12 => X"ae0010241430008c343c241030008eae001030008c343c001430008eae240014",
INIT_13 => X"00433834305854504c4844393531333742464a4e52565a0a0000000000002410",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"a9a8a7a6a5a4a3a2a1bd44e00200000062034202a560a4a0bd1d8404a5059c1c",
INIT_01 => X"a9a8a7a6a5a4a3a2a1a5a086c6c5c406bb00bb00ba5a1abfb9b8afaeadacabaa",
INIT_02 => X"9d9c9e979695949392919084e0029b401bbd60bb60bbbabfb9b8afaeadacabaa",
INIT_03 => X"6242030040008200e000c4e0000085a2e09f9d9c9e979695949392919002e09f",
INIT_04 => X"11100044508020a000b0b1b2bfbdbde000bf8400040000bfbd00e00040008284",
INIT_05 => X"424202c0e00040c543c686e30040420002e707080800a0bde0b0b1b2bf205040",
INIT_06 => X"44e002004042006263038440420042420242e042420240420062630302404200",
INIT_07 => X"86a5a2004000a200e000620042a74387e68740e6e7006000620042a7438700c0",
INIT_08 => X"86c0a000c0e00040e5e743424200064062004387e0a000c0e04086c64000a262",
INIT_09 => X"008220a0bfbdc0e00040e54342024606e74387e0a000e0e00040c5434207c643",
INIT_0A => X"e7aca5600a0b0c00400062000020854000824240008222428422004042420840",
INIT_0B => X"020222450022a5a54000e20040c2606242c2c300e60800004a000800004b0082",
INIT_0C => X"86c0804902a000004042c2a0bde000bfa50084000000000002000000a5008402",
INIT_0D => X"e2e3a20040a7e7e008e7e20261e780e20842496b008600000006008101c10107",
INIT_0E => X"e0e040a743c1c6e7a7636863c383c94802090607a202a20200e00040a7a5e7a3",
INIT_0F => X"14151010de1e52121640420200b0b1b2b3b4b5b6b7bebfbd60e0628004820080",
INIT_10 => X"0082004042008200400065a0c000156203c2004202444202420231e073e01794",
INIT_11 => X"764042002200404200c2a5444500820040a264c606004042000242e463034443",
INIT_12 => X"1500000240420062630302404200221500404200626303004042002242026540",
INIT_13 => X"00443935315955514d494541363232364145494d5155590d0000000000000200",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000ff0000200000010020000000ff18000b000c000a008900",
INIT_01 => X"00000000000000000000f8200000002000d800d800ff70000000000000000000",
INIT_02 => X"0000000000000000000000600060600000000000000000000000000000000000",
INIT_03 => X"0000200000000000000000002010000000000000000000000000000000000000",
INIT_04 => X"10000000109000888000000000ff00000000090000000000ff000000ff000000",
INIT_05 => X"000020100000ff100000100000000000000020002030000000000000001010ff",
INIT_06 => X"00002000ff0000000020000000000000200000000020ff000000002020000000",
INIT_07 => X"180000300000000000101000001000100010ff10000000000000001000103800",
INIT_08 => X"10380030100000ff100030ffff001100000000103000381000001000ff000000",
INIT_09 => X"2800004800ff100000ff1030ff101010000010300038100000ff1038ff100000",
INIT_0A => X"000000380000000000000010000018000000ffff000000000000000000ff0000",
INIT_0B => X"000000100000ff00ff0000000000001800ff0000000000000000000000000000",
INIT_0C => X"00001809000000400000ff3800000000ff0100000000010000000000ff010000",
INIT_0D => X"000000000010ff00000000000000ff000000101058000000200000008000ff00",
INIT_0E => X"1000001000ffff0010001800181818090000000000000000100000ff1000ff00",
INIT_0F => X"2000002000300020100000300000000000000000000000ff100018ff20001800",
INIT_10 => X"00800000000000000000101800280000300001cca80000200000008800982000",
INIT_11 => X"100000000000ff00000000001000800000100000200000000000000000120010",
INIT_12 => X"0000ff00ff000000002000ff0000000000ff00000000200000000000000010ff",
INIT_13 => X"00454136325a56524e4a4642373331353944484c5054580000000000000000ff",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"302c2824201c181410984408001200e84c004c0004fd2a00f80010000800ed01",
INIT_01 => X"302c2824201c181410000924504c400060125c1058fc0054504c4844403c3834",
INIT_02 => X"2824201c1814100c080400000800000801681360115c5854504c4844403c3834",
INIT_03 => X"00ff000009000000080c000810121900082c2824201c1814100c08040000082c",
INIT_04 => X"2a01cf0021250825251014181ce018080010a07900007910e8000800fa000001",
INIT_05 => X"000800250800f52a00012100000808000004000800251120081014181c2521fb",
INIT_06 => X"00080000fc0100000800ff080100000800ff08000400fc080000080000080800",
INIT_07 => X"210100250900000008252302002100210621f52a01000500070000210021250e",
INIT_08 => X"21250a25250800f32a0121c9d00200033a000021250f252508002101f9000000",
INIT_09 => X"2500002510e8250800f62a21d0402180010021250c25250800f82a21d0400100",
INIT_0A => X"010c012562780100220000253c0021040000d0f600000001010000090ad06412",
INIT_0B => X"067800210000ff01e60000000647082507c6300000620b000300781000030001",
INIT_0C => X"1a0225a400002c250323fe2518080010fe1c020004002a000500000bfe090262",
INIT_0D => X"000000000a2bff000101002d0401eb000123212312180000120d00020004ff0d",
INIT_0E => X"2508002100f6fc01210021ff062404ec000f1c0201780030250800f82b01ff00",
INIT_0F => X"0004d8000400600000000800001014181c2024282c3034c8250821fd43012505",
INIT_10 => X"00130009010000000e002a252e2500000000e0400000700000997425d4250008",
INIT_11 => X"2a2010000000f3020000010021001300060000d8000011020000000001830021",
INIT_12 => X"0000a999fc100000740099b21000000000fc1000007400000810000000cc2ad5",
INIT_13 => X"00464237330057534f4b4743383430343843474b4f535700000000000000cce2",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
