-------------------------------------------------------------------------------
-- Inferred BlockRAM with Initial Values
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Ram_Program is
  generic (
    N : integer := 4;                -- Width in bytes
    M : integer := 13);               -- Address width

  port (
    clk  : in  std_logic;
    wbe   : in  std_logic_vector(N-1 downto 0)   := (others => '0');
    addr : in  std_logic_vector(M-1 downto 0)   := (others => '0');
    din  : in  std_logic_vector(N*8-1 downto 0) := (others => '0');
    dout : out std_logic_vector(N*8-1 downto 0)
    );

end Ram_Program;

architecture logic of Ram_Program is

  type mem_file is array(0 to (2**M)-1) of std_logic_vector(N*8-1 downto 0);
  
  signal ram : mem_file := (
    -- Insert initial values below here, eg,
    -- 0 => X"0000",
    -- 1 => X"0001",
    -- <INIT_DATA>
0 => X"3C1C0001",1 => X"279CA274",2 => X"3C050000",3 => X"24A522B0",
4 => X"3C040000",5 => X"248423C0",6 => X"341D8000",7 => X"ACA00000",
8 => X"00A4182A",9 => X"1460FFFD",10 => X"24A50004",11 => X"3C020000",
12 => X"2442005C",13 => X"3C032000",14 => X"AC62004C",15 => X"0C000741",
16 => X"00000000",17 => X"08000011",18 => X"00000000",19 => X"3C020000",
20 => X"244223C0",21 => X"03E00008",22 => X"00000000",23 => X"3C022000",
24 => X"03E00008",25 => X"AC440044",26 => X"40026000",27 => X"03E00008",
28 => X"40846000",29 => X"00000000",30 => X"00000000",31 => X"00000000",
32 => X"23BDFF98",33 => X"AFA10010",34 => X"AFA20014",35 => X"AFA30018",
36 => X"AFA4001C",37 => X"AFA50020",38 => X"AFA60024",39 => X"AFA70028",
40 => X"AFA8002C",41 => X"AFA90030",42 => X"AFAA0034",43 => X"AFAB0038",
44 => X"AFAC003C",45 => X"AFAD0040",46 => X"AFAE0044",47 => X"AFAF0048",
48 => X"AFB8004C",49 => X"AFB90050",50 => X"AFBF0054",51 => X"401A7000",
52 => X"235AFFFC",53 => X"AFBA0058",54 => X"0000D810",55 => X"AFBB005C",
56 => X"0000D812",57 => X"AFBB0060",58 => X"3C062000",59 => X"8CC40040",
60 => X"8CC5004C",61 => X"8CC60050",62 => X"00862024",63 => X"00A0F809",
64 => X"23A50000",65 => X"8FA10010",66 => X"8FA20014",67 => X"8FA30018",
68 => X"8FA4001C",69 => X"8FA50020",70 => X"8FA60024",71 => X"8FA70028",
72 => X"8FA8002C",73 => X"8FA90030",74 => X"8FAA0034",75 => X"8FAB0038",
76 => X"8FAC003C",77 => X"8FAD0040",78 => X"8FAE0044",79 => X"8FAF0048",
80 => X"8FB8004C",81 => X"8FB90050",82 => X"8FBF0054",83 => X"8FBA0058",
84 => X"8FBB005C",85 => X"03600011",86 => X"8FBB0060",87 => X"03600013",
88 => X"23BD0068",89 => X"341B0001",90 => X"03400008",91 => X"409B6000",
92 => X"AC900000",93 => X"AC910004",94 => X"AC920008",95 => X"AC93000C",
96 => X"AC940010",97 => X"AC950014",98 => X"AC960018",99 => X"AC97001C",
100 => X"AC9E0020",101 => X"AC9C0024",102 => X"AC9D0028",103 => X"AC9F002C",
104 => X"03E00008",105 => X"34020000",106 => X"8C900000",107 => X"8C910004",
108 => X"8C920008",109 => X"8C93000C",110 => X"8C940010",111 => X"8C950014",
112 => X"8C960018",113 => X"8C97001C",114 => X"8C9E0020",115 => X"8C9C0024",
116 => X"8C9D0028",117 => X"8C9F002C",118 => X"03E00008",119 => X"34A20000",
120 => X"00850019",121 => X"00001012",122 => X"00002010",123 => X"03E00008",
124 => X"ACC40000",125 => X"0000000C",126 => X"03E00008",127 => X"00000000",
128 => X"90820000",129 => X"00000000",130 => X"10400009",131 => X"00000000",
132 => X"3C032000",133 => X"304200FF",134 => X"AC620000",135 => X"24840001",
136 => X"90820000",137 => X"00000000",138 => X"1440FFFA",139 => X"00000000",
140 => X"03E00008",141 => X"00000000",142 => X"27BDFFE8",143 => X"AFBF0010",
144 => X"0C000080",145 => X"00000000",146 => X"3C040000",147 => X"0C000080",
148 => X"248421A0",149 => X"8FBF0010",150 => X"00000000",151 => X"03E00008",
152 => X"27BD0018",153 => X"27BDFFE0",154 => X"AFBF001C",155 => X"AFB20018",
156 => X"AFB10014",157 => X"AFB00010",158 => X"00008025",159 => X"00A08825",
160 => X"1A200008",161 => X"00809025",162 => X"02501021",163 => X"90440000",
164 => X"0C0000D6",165 => X"26100001",166 => X"0211102A",167 => X"1440FFFB",
168 => X"02501021",169 => X"02201025",170 => X"8FBF001C",171 => X"8FB20018",
172 => X"8FB10014",173 => X"8FB00010",174 => X"03E00008",175 => X"27BD0020",
176 => X"18A00011",177 => X"00003025",178 => X"3C082000",179 => X"35080008",
180 => X"3C072000",181 => X"34E70004",182 => X"8D020000",183 => X"00000000",
184 => X"30420008",185 => X"10400008",186 => X"00000000",187 => X"8CE30000",
188 => X"00861021",189 => X"24C60001",190 => X"A0430000",191 => X"00C5102A",
192 => X"1440FFF5",193 => X"00000000",194 => X"03E00008",195 => X"00C01025",
196 => X"3C022000",197 => X"34420008",198 => X"8C420000",199 => X"00000000",
200 => X"30420008",201 => X"14400008",202 => X"3C022000",203 => X"3C032000",
204 => X"34630008",205 => X"8C620000",206 => X"00000000",207 => X"30420008",
208 => X"1040FFFC",209 => X"3C022000",210 => X"34420004",211 => X"8C420000",
212 => X"03E00008",213 => X"304200FF",214 => X"3C022000",215 => X"34420008",
216 => X"8C420000",217 => X"00000000",218 => X"30420001",219 => X"10400008",
220 => X"308400FF",221 => X"3C032000",222 => X"34630008",223 => X"8C620000",
224 => X"00000000",225 => X"30420001",226 => X"1440FFFC",227 => X"00000000",
228 => X"3C022000",229 => X"03E00008",230 => X"AC440000",231 => X"18C0000E",
232 => X"00003825",233 => X"00871021",234 => X"90430000",235 => X"00A71021",
236 => X"90420000",237 => X"00000000",238 => X"14620007",239 => X"00000000",
240 => X"10600005",241 => X"00000000",242 => X"24E70001",243 => X"00E6102A",
244 => X"1440FFF5",245 => X"00871021",246 => X"10E60006",247 => X"00871021",
248 => X"90430000",249 => X"00A71021",250 => X"90420000",251 => X"10000002",
252 => X"00621023",253 => X"00001025",254 => X"03E00008",255 => X"00000000",
256 => X"90A20000",257 => X"00000000",258 => X"10400009",259 => X"00003025",
260 => X"90A20000",261 => X"24A50001",262 => X"00861821",263 => X"A0620000",
264 => X"90A20000",265 => X"00000000",266 => X"1440FFF9",267 => X"24C60001",
268 => X"00861021",269 => X"A0400000",270 => X"03E00008",271 => X"00C01025",
272 => X"00003825",273 => X"18A0000F",274 => X"00E03025",275 => X"00871021",
276 => X"90430000",277 => X"00000000",278 => X"2C62003A",279 => X"10400003",
280 => X"00061100",281 => X"10000002",282 => X"2442FFD0",283 => X"2442FFC9",
284 => X"00433021",285 => X"24E70001",286 => X"00E5102A",287 => X"1440FFF3",
288 => X"00000000",289 => X"03E00008",290 => X"00C01025",291 => X"00003025",
292 => X"18A0000A",293 => X"00C03825",294 => X"00861021",295 => X"90430000",
296 => X"24C60001",297 => X"00071040",298 => X"2442FFD0",299 => X"00433821",
300 => X"00C5102A",301 => X"1440FFF8",302 => X"00000000",303 => X"03E00008",
304 => X"00E01025",305 => X"00003825",306 => X"18A0000C",307 => X"00E03025",
308 => X"00871021",309 => X"90430000",310 => X"24E70001",311 => X"00061080",
312 => X"00461021",313 => X"00021040",314 => X"2442FFD0",315 => X"00433021",
316 => X"00E5102A",317 => X"1440FFF6",318 => X"00000000",319 => X"03E00008",
320 => X"00C01025",321 => X"27BDFFE8",322 => X"AFBF0010",323 => X"00A04825",
324 => X"AD200000",325 => X"90820000",326 => X"00002825",327 => X"10400012",
328 => X"24080064",329 => X"2442FFD0",330 => X"2C42000A",331 => X"14400009",
332 => X"00000000",333 => X"8D220000",334 => X"24840001",335 => X"24420001",
336 => X"AD220000",337 => X"90820000",338 => X"00000000",339 => X"1440FFF6",
340 => X"2442FFD0",341 => X"90820000",342 => X"00000000",343 => X"14400004",
344 => X"00851821",345 => X"AD200000",346 => X"1000003C",347 => X"00001025",
348 => X"90620000",349 => X"00000000",350 => X"10400022",351 => X"00000000",
352 => X"240C0001",353 => X"240B0078",354 => X"240A0062",355 => X"00603825",
356 => X"24A50001",357 => X"14AC000C",358 => X"24E70001",359 => X"90820001",
360 => X"00000000",361 => X"144B0003",362 => X"00000000",363 => X"10000010",
364 => X"24080078",365 => X"00000000",366 => X"144A0003",367 => X"00000000",
368 => X"1000000B",369 => X"24080062",370 => X"90E60000",371 => X"00000000",
372 => X"2CC30030",373 => X"24C2FFC6",374 => X"2C420007",375 => X"00621825",
376 => X"14600008",377 => X"2CC20047",378 => X"10400006",379 => X"00000000",
380 => X"90E20000",381 => X"00000000",382 => X"1440FFE6",383 => X"24A50001",
384 => X"24A5FFFF",385 => X"8D220000",386 => X"00000000",387 => X"00451021",
388 => X"AD220000",389 => X"24020078",390 => X"15020006",391 => X"24020062",
392 => X"24840002",393 => X"0C000110",394 => X"24A5FFFE",395 => X"1000000B",
396 => X"00000000",397 => X"00000000",398 => X"11020005",399 => X"00000000",
400 => X"0C000131",401 => X"00000000",402 => X"10000004",403 => X"00000000",
404 => X"24840002",405 => X"0C000123",406 => X"24A5FFFE",407 => X"8FBF0010",
408 => X"00000000",409 => X"03E00008",410 => X"27BD0018",411 => X"00A03825",
412 => X"24C2FFFE",413 => X"2C420023",414 => X"14400003",415 => X"00004025",
416 => X"1000002C",417 => X"A0A00000",418 => X"3C020000",419 => X"244921A4",
420 => X"00801825",421 => X"14C00002",422 => X"0086001A",423 => X"0007000D",
424 => X"2401FFFF",425 => X"14C10004",426 => X"3C018000",427 => X"14810002",
428 => X"00000000",429 => X"0006000D",430 => X"00002012",431 => X"00000000",
432 => X"00000000",433 => X"00860018",434 => X"00005812",435 => X"006B1023",
436 => X"00491021",437 => X"90420023",438 => X"25080001",439 => X"A0E20000",
440 => X"1480FFEB",441 => X"24E70001",442 => X"04610004",443 => X"2402002D",
444 => X"A0E20000",445 => X"24E70001",446 => X"25080001",447 => X"A0E00000",
448 => X"24E7FFFF",449 => X"00A7102B",450 => X"1040000A",451 => X"00000000",
452 => X"90A20000",453 => X"90E30000",454 => X"A0E20000",455 => X"A0A30000",
456 => X"24E7FFFF",457 => X"24A50001",458 => X"00A7102B",459 => X"1440FFF8",
460 => X"00000000",461 => X"03E00008",462 => X"01001025",463 => X"24020030",
464 => X"A0A20000",465 => X"24020078",466 => X"A0A20001",467 => X"24070002",
468 => X"2406001C",469 => X"2409000F",470 => X"3C020000",471 => X"244821EC",
472 => X"00C91804",473 => X"00831824",474 => X"00C31806",475 => X"306300FF",
476 => X"00681821",477 => X"90630000",478 => X"00A71021",479 => X"24E70001",
480 => X"24C6FFFC",481 => X"04C1FFF6",482 => X"A0430000",483 => X"00A71021",
484 => X"A0400000",485 => X"03E00008",486 => X"00E01025",487 => X"18C00016",
488 => X"00003825",489 => X"3C020000",490 => X"244921EC",491 => X"24A80001",
492 => X"00871821",493 => X"90620000",494 => X"00000000",495 => X"00021102",
496 => X"00491021",497 => X"90420000",498 => X"00000000",499 => X"A0A20000",
500 => X"90620000",501 => X"24E70001",502 => X"3042000F",503 => X"00491021",
504 => X"90420000",505 => X"24A50002",506 => X"A1020000",507 => X"00E6102A",
508 => X"1440FFEF",509 => X"25080002",510 => X"03E00008",511 => X"00000000",
512 => X"3C022000",513 => X"34420044",514 => X"AC440000",515 => X"8F828024",
516 => X"3C032000",517 => X"34630060",518 => X"24420001",519 => X"AF828024",
520 => X"03E00008",521 => X"AC620000",522 => X"27BDFFE8",523 => X"AFBF0010",
524 => X"3C022000",525 => X"34420060",526 => X"AC440000",527 => X"28822711",
528 => X"14400006",529 => X"00000000",530 => X"3C040000",531 => X"0C000080",
532 => X"24842200",533 => X"10000003",534 => X"00000000",535 => X"0C00020A",
536 => X"24840001",537 => X"8FBF0010",538 => X"00000000",539 => X"03E00008",
540 => X"27BD0018",541 => X"27BDFFE8",542 => X"AFBF0010",543 => X"0C000013",
544 => X"00000000",545 => X"AF82803C",546 => X"00402825",547 => X"3C042000",
548 => X"34840060",549 => X"00051E03",550 => X"AC830000",551 => X"00051C03",
552 => X"AC830000",553 => X"00051A03",554 => X"AC830000",555 => X"AC850000",
556 => X"24050063",557 => X"2442018C",558 => X"AC450000",559 => X"24A5FFFF",
560 => X"04A1FFFD",561 => X"2442FFFC",562 => X"00002825",563 => X"3C032000",
564 => X"34630060",565 => X"AC650000",566 => X"24A50001",567 => X"28A20064",
568 => X"1440FFFC",569 => X"00000000",570 => X"8FBF0010",571 => X"00000000",
572 => X"03E00008",573 => X"27BD0018",574 => X"8C820010",575 => X"00000000",
576 => X"ACA20004",577 => X"8C82000C",578 => X"00000000",579 => X"ACA20000",
580 => X"90820009",581 => X"03E00008",582 => X"A0A20008",583 => X"8C820004",
584 => X"00000000",585 => X"ACA20004",586 => X"8C820000",587 => X"00000000",
588 => X"ACA20000",589 => X"90820008",590 => X"03E00008",591 => X"A0A20008",
592 => X"8CA30000",593 => X"00000000",594 => X"10600005",595 => X"00000000",
596 => X"8C820000",597 => X"00000000",598 => X"14620012",599 => X"00001025",
600 => X"8CA30004",601 => X"00000000",602 => X"10600005",603 => X"00000000",
604 => X"8C820004",605 => X"00000000",606 => X"1462000A",607 => X"00001025",
608 => X"90A50008",609 => X"00000000",610 => X"10A00006",611 => X"24020001",
612 => X"90830008",613 => X"00000000",614 => X"14A30002",615 => X"00001025",
616 => X"24020001",617 => X"03E00008",618 => X"00000000",619 => X"27BDFFD8",
620 => X"AFBF0024",621 => X"AFB20020",622 => X"AFB1001C",623 => X"AFB00018",
624 => X"00808825",625 => X"0C000141",626 => X"27A50010",627 => X"8FB00010",
628 => X"00409025",629 => X"27A50010",630 => X"0C000141",631 => X"02302021",
632 => X"00121A00",633 => X"00629021",634 => X"8FA20010",635 => X"27A50010",
636 => X"02028021",637 => X"0C000141",638 => X"02302021",639 => X"00121A00",
640 => X"00629021",641 => X"8FA20010",642 => X"27A50010",643 => X"02028021",
644 => X"0C000141",645 => X"02302021",646 => X"8FBF0024",647 => X"00121A00",
648 => X"8FB20020",649 => X"8FB1001C",650 => X"8FB00018",651 => X"00621021",
652 => X"03E00008",653 => X"27BD0028",654 => X"27BDFFE0",655 => X"AFBF0018",
656 => X"AFB10014",657 => X"AFB00010",658 => X"AFA40020",659 => X"27A40020",
660 => X"00A08025",661 => X"0C0001E7",662 => X"24060001",663 => X"2411002E",
664 => X"A2110002",665 => X"27A40021",666 => X"26050003",667 => X"0C0001E7",
668 => X"24060001",669 => X"A2110005",670 => X"27A40022",671 => X"26050006",
672 => X"0C0001E7",673 => X"24060001",674 => X"A2110008",675 => X"27A40023",
676 => X"26050009",677 => X"0C0001E7",678 => X"24060001",679 => X"8FBF0018",
680 => X"8FB10014",681 => X"8FB00010",682 => X"03E00008",683 => X"27BD0020",
684 => X"27BDFFC8",685 => X"AFBF0030",686 => X"AFB5002C",687 => X"AFB40028",
688 => X"AFB30024",689 => X"AFB20020",690 => X"AFB1001C",691 => X"AFB00018",
692 => X"00808825",693 => X"3C040000",694 => X"2484220C",695 => X"0C000099",
696 => X"24050002",697 => X"3C020000",698 => X"245022C0",699 => X"8E220020",
700 => X"27A40010",701 => X"02002825",702 => X"24060004",703 => X"0C0001E7",
704 => X"AFA20010",705 => X"02002025",706 => X"0C000099",707 => X"24050008",
708 => X"0C0000D6",709 => X"2404003B",710 => X"8FA30010",711 => X"8F828040",
712 => X"00000000",713 => X"14620053",714 => X"02002825",715 => X"8E24002C",
716 => X"0C00028E",717 => X"AFA40010",718 => X"02002025",719 => X"0C000099",
720 => X"2405000B",721 => X"0C0000D6",722 => X"2404003B",723 => X"93828030",
724 => X"00000000",725 => X"14400004",726 => X"00000000",727 => X"8FA20010",
728 => X"00000000",729 => X"AF82802C",730 => X"8E240030",731 => X"02002825",
732 => X"0C00028E",733 => X"AFA40010",734 => X"02002025",735 => X"0C000099",
736 => X"2405000B",737 => X"0C0000D6",738 => X"2404003B",739 => X"93828030",
740 => X"00000000",741 => X"14400004",742 => X"00000000",743 => X"8FA20010",
744 => X"00000000",745 => X"AF828034",746 => X"2631010C",747 => X"00009025",
748 => X"241500FF",749 => X"24140001",750 => X"02009825",751 => X"92230000",
752 => X"00000000",753 => X"1075002B",754 => X"00000000",755 => X"92300001",
756 => X"00000000",757 => X"2E020020",758 => X"10400026",759 => X"38630033",
760 => X"2C630001",761 => X"3A020004",762 => X"2C420001",763 => X"00621824",
764 => X"10600010",765 => X"00000000",766 => X"93828030",767 => X"00000000",
768 => X"1454000C",769 => X"00000000",770 => X"92220002",771 => X"92230003",
772 => X"92240004",773 => X"92250005",774 => X"00021600",775 => X"00031C00",
776 => X"00431021",777 => X"00042200",778 => X"00441021",779 => X"00451021",
780 => X"AF828028",781 => X"02202025",782 => X"02602825",783 => X"0C0001E7",
784 => X"26060002",785 => X"02602025",786 => X"00102840",787 => X"0C000099",
788 => X"24A50004",789 => X"0C0000D6",790 => X"2404003B",791 => X"02301021",
792 => X"24510002",793 => X"26520001",794 => X"2A42000A",795 => X"1440FFD3",
796 => X"00000000",797 => X"8FBF0030",798 => X"8FB5002C",799 => X"8FB40028",
800 => X"8FB30024",801 => X"8FB20020",802 => X"8FB1001C",803 => X"8FB00018",
804 => X"03E00008",805 => X"27BD0038",806 => X"27BDFFE0",807 => X"AFBF0018",
808 => X"AFB10014",809 => X"AFB00010",810 => X"00808025",811 => X"3C040000",
812 => X"24842210",813 => X"00A08825",814 => X"0C000099",815 => X"24050002",
816 => X"26040014",817 => X"3C100000",818 => X"261022C0",819 => X"02002825",
820 => X"0C0001E7",821 => X"24060002",822 => X"02002025",823 => X"0C000099",
824 => X"24050004",825 => X"0C0000D6",826 => X"2404003B",827 => X"8F838038",
828 => X"24020003",829 => X"10620010",830 => X"00000000",831 => X"8F828038",
832 => X"02202025",833 => X"3C100000",834 => X"24420001",835 => X"AF828038",
836 => X"8F858038",837 => X"26102340",838 => X"00052940",839 => X"0C000247",
840 => X"00B02821",841 => X"8F828038",842 => X"00000000",843 => X"00021140",
844 => X"00501021",845 => X"AC40001C",846 => X"8FBF0018",847 => X"8FB10014",
848 => X"8FB00010",849 => X"03E00008",850 => X"27BD0020",851 => X"27BDFFE8",
852 => X"AFBF0014",853 => X"AFB00010",854 => X"00808025",855 => X"0C0000D6",
856 => X"24040054",857 => X"26040014",858 => X"3C100000",859 => X"261022C0",
860 => X"02002825",861 => X"0C0001E7",862 => X"24060002",863 => X"02002025",
864 => X"0C000099",865 => X"24050004",866 => X"0C0000D6",867 => X"2404003B",
868 => X"8FBF0014",869 => X"8FB00010",870 => X"03E00008",871 => X"27BD0018",
872 => X"27BDFFD8",873 => X"AFBF0020",874 => X"AFB1001C",875 => X"AFB00018",
876 => X"00808825",877 => X"96220014",878 => X"96230016",879 => X"3C040000",
880 => X"24842214",881 => X"24050002",882 => X"A7A20010",883 => X"0C000099",
884 => X"A7A30012",885 => X"27A40010",886 => X"3C100000",887 => X"261022C0",
888 => X"02002825",889 => X"0C0001E7",890 => X"24060002",891 => X"02002025",
892 => X"0C000099",893 => X"24050004",894 => X"0C0000D6",895 => X"2404003B",
896 => X"27A40012",897 => X"02002825",898 => X"0C0001E7",899 => X"24060002",
900 => X"02002025",901 => X"0C000099",902 => X"24050004",903 => X"0C0000D6",
904 => X"2404003B",905 => X"97A30012",906 => X"24020044",907 => X"14620003",
908 => X"00000000",909 => X"0C0002AC",910 => X"02202025",911 => X"8FBF0020",
912 => X"8FB1001C",913 => X"8FB00018",914 => X"03E00008",915 => X"27BD0028",
916 => X"27BDFFE8",917 => X"AFBF0014",918 => X"AFB00010",919 => X"00808025",
920 => X"3C040000",921 => X"24842218",922 => X"0C000099",923 => X"24050002",
924 => X"26040014",925 => X"3C100000",926 => X"261022C0",927 => X"02002825",
928 => X"0C0001E7",929 => X"24060002",930 => X"02002025",931 => X"0C000099",
932 => X"24050004",933 => X"0C0000D6",934 => X"2404003B",935 => X"8FBF0014",
936 => X"8FB00010",937 => X"03E00008",938 => X"27BD0018",939 => X"27BDFFE8",
940 => X"AFBF0014",941 => X"AFB00010",942 => X"00A08025",943 => X"3C040000",
944 => X"2484221C",945 => X"0C000099",946 => X"24050002",947 => X"8F838038",
948 => X"24020003",949 => X"10620023",950 => X"00000000",951 => X"8F828038",
952 => X"3C052001",953 => X"34A55034",954 => X"3C062001",955 => X"34C65038",
956 => X"3C072001",957 => X"34E7503C",958 => X"3C040000",959 => X"24842340",
960 => X"24030001",961 => X"02052826",962 => X"02063026",963 => X"24420001",
964 => X"AF828038",965 => X"8F828038",966 => X"02073826",967 => X"00021140",
968 => X"00441021",969 => X"AC43001C",970 => X"8F828038",971 => X"8CA30000",
972 => X"00021140",973 => X"00441021",974 => X"AC43000C",975 => X"8F828038",
976 => X"8CC30000",977 => X"00021140",978 => X"00441021",979 => X"AC430010",
980 => X"8F828038",981 => X"8CE30000",982 => X"00021140",983 => X"00441021",
984 => X"AC430014",985 => X"8FBF0014",986 => X"8FB00010",987 => X"03E00008",
988 => X"27BD0018",989 => X"27BDFFB8",990 => X"AFBF0044",991 => X"AFBE0040",
992 => X"AFB7003C",993 => X"AFB60038",994 => X"AFB50034",995 => X"AFB40030",
996 => X"AFB3002C",997 => X"AFB20028",998 => X"AFB10024",999 => X"AFB00020",
1000 => X"AFA40048",1001 => X"00008825",1002 => X"3C132001",1003 => X"36735020",
1004 => X"3C020000",1005 => X"245222C0",1006 => X"241E003B",1007 => X"3C170000",
1008 => X"24160011",1009 => X"24150001",1010 => X"24140006",1011 => X"02331026",
1012 => X"8C420000",1013 => X"00000000",1014 => X"3042FFFF",1015 => X"10400082",
1016 => X"3C022001",1017 => X"34425030",1018 => X"02221026",1019 => X"8C420000",
1020 => X"3C032001",1021 => X"34634000",1022 => X"02238026",1023 => X"3043FFFF",
1024 => X"24020800",1025 => X"1462002D",1026 => X"00602025",1027 => X"02002025",
1028 => X"0C00023E",1029 => X"27A50010",1030 => X"3C070000",1031 => X"24E42220",
1032 => X"0C000099",1033 => X"24050003",1034 => X"8FA40010",1035 => X"A25E000B",
1036 => X"0C00028E",1037 => X"02402825",1038 => X"02402025",1039 => X"0C000099",
1040 => X"2405000C",1041 => X"8FA40014",1042 => X"0C00028E",1043 => X"02402825",
1044 => X"02402025",1045 => X"0C000099",1046 => X"2405000C",1047 => X"27A40018",
1048 => X"02402825",1049 => X"0C0001E7",1050 => X"24060001",1051 => X"02402025",
1052 => X"0C000099",1053 => X"24050002",1054 => X"0C0000D6",1055 => X"2404003B",
1056 => X"27A40010",1057 => X"0C000250",1058 => X"26E52278",1059 => X"10400057",
1060 => X"02331026",1061 => X"93A20018",1062 => X"00000000",1063 => X"10560037",
1064 => X"02002025",1065 => X"1055003C",1066 => X"00000000",1067 => X"10540040",
1068 => X"00000000",1069 => X"10000042",1070 => X"00000000",1071 => X"24020806",
1072 => X"10620046",1073 => X"2C820600",1074 => X"10400047",1075 => X"3C02F000",
1076 => X"8E040000",1077 => X"3C034000",1078 => X"00821024",1079 => X"1443003C",
1080 => X"3C020001",1081 => X"02002025",1082 => X"0C00023E",1083 => X"27A50010",
1084 => X"3C070000",1085 => X"24E42220",1086 => X"0C000099",1087 => X"24050003",
1088 => X"8FA40010",1089 => X"A25E000B",1090 => X"0C00028E",1091 => X"02402825",
1092 => X"02402025",1093 => X"0C000099",1094 => X"2405000C",1095 => X"8FA40014",
1096 => X"0C00028E",1097 => X"02402825",1098 => X"02402025",1099 => X"0C000099",
1100 => X"2405000C",1101 => X"27A40018",1102 => X"02402825",1103 => X"0C0001E7",
1104 => X"24060001",1105 => X"02402025",1106 => X"0C000099",1107 => X"24050002",
1108 => X"0C0000D6",1109 => X"2404003B",1110 => X"27A40010",1111 => X"0C000250",
1112 => X"26E52278",1113 => X"10400021",1114 => X"02331026",1115 => X"93A20018",
1116 => X"00000000",1117 => X"14560005",1118 => X"02002025",1119 => X"0C000368",
1120 => X"27A50010",1121 => X"10000019",1122 => X"02331026",1123 => X"00000000",
1124 => X"14550005",1125 => X"00000000",1126 => X"0C000326",1127 => X"27A50010",
1128 => X"10000012",1129 => X"02331026",1130 => X"14540005",1131 => X"02002025",
1132 => X"0C000353",1133 => X"27A50010",1134 => X"1000000C",1135 => X"02331026",
1136 => X"0C000394",1137 => X"27A50010",1138 => X"10000008",1139 => X"02331026",
1140 => X"34420800",1141 => X"14820005",1142 => X"02331026",1143 => X"02002025",
1144 => X"0C0003AB",1145 => X"02202825",1146 => X"02331026",1147 => X"AC400000",
1148 => X"26310800",1149 => X"2E220801",1150 => X"1440FF75",1151 => X"02331026",
1152 => X"8F828018",1153 => X"8FA70048",1154 => X"00000000",1155 => X"AC470000",
1156 => X"8FBF0044",1157 => X"8FBE0040",1158 => X"8FB7003C",1159 => X"8FB60038",
1160 => X"8FB50034",1161 => X"8FB40030",1162 => X"8FB3002C",1163 => X"8FB20028",
1164 => X"8FB10024",1165 => X"8FB00020",1166 => X"03E00008",1167 => X"27BD0048",
1168 => X"27BDFFE8",1169 => X"AFBF0010",1170 => X"3C022001",1171 => X"34420024",
1172 => X"3084FFFF",1173 => X"AC440000",1174 => X"3C022001",1175 => X"34420028",
1176 => X"30A5FFFF",1177 => X"AC450000",1178 => X"3C022001",1179 => X"3442002C",
1180 => X"30C6FFFF",1181 => X"AC460000",1182 => X"3C022001",1183 => X"34425020",
1184 => X"AC400000",1185 => X"3C022001",1186 => X"34425820",1187 => X"AC400000",
1188 => X"8F83801C",1189 => X"3C020000",1190 => X"24420F74",1191 => X"AC620000",
1192 => X"8F838020",1193 => X"24020004",1194 => X"AC620000",1195 => X"8F828014",
1196 => X"24040001",1197 => X"0C00001A",1198 => X"AC400000",1199 => X"8FBF0010",
1200 => X"00000000",1201 => X"03E00008",1202 => X"27BD0018",1203 => X"00001825",
1204 => X"30A5FFFF",1205 => X"10A00008",1206 => X"00603025",1207 => X"94820000",
1208 => X"24630002",1209 => X"3063FFFF",1210 => X"00C23021",1211 => X"0065102B",
1212 => X"1440FFFA",1213 => X"24840002",1214 => X"30C3FFFF",1215 => X"00061402",
1216 => X"00623021",1217 => X"00061027",1218 => X"03E00008",1219 => X"3042FFFF",
1220 => X"3C022001",1221 => X"34423024",1222 => X"3084FFFF",1223 => X"AC440000",
1224 => X"3C022001",1225 => X"34423028",1226 => X"30A5FFFF",1227 => X"AC450000",
1228 => X"3C022001",1229 => X"3442302C",1230 => X"30C6FFFF",1231 => X"03E00008",
1232 => X"AC460000",1233 => X"27BDFFE8",1234 => X"AFBF0014",1235 => X"AFB00010",
1236 => X"24024500",1237 => X"3C012001",1238 => X"A4222000",1239 => X"3C012001",
1240 => X"A4242002",1241 => X"3C026DF3",1242 => X"3C012001",1243 => X"AC222004",
1244 => X"30A580FF",1245 => X"34A58000",1246 => X"3C012001",1247 => X"A4252008",
1248 => X"3C102001",1249 => X"3610200A",1250 => X"A6000000",1251 => X"3C012001",
1252 => X"AC26200C",1253 => X"3C012001",1254 => X"AC272010",1255 => X"3C042001",
1256 => X"34842000",1257 => X"0C0004B3",1258 => X"24050014",1259 => X"A6020000",
1260 => X"8FBF0014",1261 => X"8FB00010",1262 => X"03E00008",1263 => X"27BD0018",
1264 => X"27BDFFE0",1265 => X"AFBF0018",1266 => X"AFB10014",1267 => X"AFB00010",
1268 => X"00801825",1269 => X"00C08825",1270 => X"3224FFFF",1271 => X"00A01025",
1272 => X"24050001",1273 => X"00E08025",1274 => X"3210FFFF",1275 => X"00603025",
1276 => X"0C0004D1",1277 => X"00403825",1278 => X"24020800",1279 => X"3C012001",
1280 => X"A4222014",1281 => X"3C012001",1282 => X"A4202016",1283 => X"24020001",
1284 => X"3C012001",1285 => X"A4222018",1286 => X"3C012001",1287 => X"A430201A",
1288 => X"3C042001",1289 => X"3484201C",1290 => X"2625FFE4",1291 => X"18A00008",
1292 => X"00001825",1293 => X"3062000F",1294 => X"24420061",1295 => X"A0820000",
1296 => X"24630001",1297 => X"0065102A",1298 => X"1440FFFA",1299 => X"24840001",
1300 => X"3C042001",1301 => X"34842014",1302 => X"2625FFEC",1303 => X"0C0004B3",
1304 => X"30A5FFFF",1305 => X"8FBF0018",1306 => X"8FB10014",1307 => X"8FB00010",
1308 => X"3C012001",1309 => X"A4222016",1310 => X"03E00008",1311 => X"27BD0020",
1312 => X"27BDFFD8",1313 => X"AFB20018",1314 => X"8FB20038",1315 => X"AFBF0024",
1316 => X"AFB40020",1317 => X"AFB3001C",1318 => X"AFB10014",1319 => X"AFB00010",
1320 => X"3C132001",1321 => X"36732014",1322 => X"00801025",1323 => X"00A01825",
1324 => X"00C08025",1325 => X"00E08825",1326 => X"3210FFFF",1327 => X"3231FFFF",
1328 => X"24050011",1329 => X"00403025",1330 => X"00603825",1331 => X"2654001C",
1332 => X"0C0004D1",1333 => X"3284FFFF",1334 => X"A6700000",1335 => X"A6710002",
1336 => X"26520008",1337 => X"A6720004",1338 => X"A6600006",1339 => X"8FBF0024",
1340 => X"02801025",1341 => X"8FB40020",1342 => X"8FB3001C",1343 => X"8FB20018",
1344 => X"8FB10014",1345 => X"8FB00010",1346 => X"03E00008",1347 => X"27BD0028",
1348 => X"27BDFFE0",1349 => X"AFBF001C",1350 => X"AFB00018",1351 => X"00808025",
1352 => X"3404FFFF",1353 => X"00802825",1354 => X"0C0004C4",1355 => X"00803025",
1356 => X"3C052001",1357 => X"34A5201C",1358 => X"3C020101",1359 => X"34420600",
1360 => X"ACA20000",1361 => X"3C012001",1362 => X"AC302020",1363 => X"3C012001",
1364 => X"AC202024",1365 => X"3C012001",1366 => X"AC202028",1367 => X"3C012001",
1368 => X"AC20202C",1369 => X"3C012001",1370 => X"AC202030",1371 => X"3C012001",
1372 => X"AC202034",1373 => X"2402020A",1374 => X"3C012001",1375 => X"A4222038",
1376 => X"24023544",1377 => X"3C012001",1378 => X"A422203A",1379 => X"24025441",
1380 => X"3C012001",1381 => X"A422203C",1382 => X"24030022",1383 => X"240400C9",
1384 => X"00A31021",1385 => X"A0400000",1386 => X"2484FFFF",1387 => X"0481FFFC",
1388 => X"24630001",1389 => X"3C026382",1390 => X"34425363",1391 => X"ACA200EC",
1392 => X"24023501",1393 => X"A4A200F0",1394 => X"24020001",1395 => X"A0A200F2",
1396 => X"240200FF",1397 => X"A0A200F3",1398 => X"240300F4",1399 => X"AFA30010",
1400 => X"00002025",1401 => X"2405FFFF",1402 => X"24060044",1403 => X"0C000520",
1404 => X"24070043",1405 => X"8FBF001C",1406 => X"8FB00018",1407 => X"03E00008",
1408 => X"27BD0020",1409 => X"8F838034",1410 => X"3C023501",1411 => X"34420300",
1412 => X"3C012001",1413 => X"AC22210C",1414 => X"24023204",1415 => X"3C012001",
1416 => X"A4222110",1417 => X"240200FF",1418 => X"3C012001",1419 => X"A0222116",
1420 => X"27BDFFE0",1421 => X"240200FB",1422 => X"AFA20010",1423 => X"8F82802C",
1424 => X"AFBF0018",1425 => X"00002025",1426 => X"2405FFFF",1427 => X"24060044",
1428 => X"24070043",1429 => X"3C012001",1430 => X"AC232030",1431 => X"8F83802C",
1432 => X"00021402",1433 => X"3C012001",1434 => X"A4222112",1435 => X"3C012001",
1436 => X"0C000520",1437 => X"A4232114",1438 => X"8FBF0018",1439 => X"00000000",
1440 => X"03E00008",1441 => X"27BD0020",1442 => X"27BDFFD8",1443 => X"AFBF0024",
1444 => X"AFB40020",1445 => X"AFB3001C",1446 => X"AFB20018",1447 => X"AFB10014",
1448 => X"AFB00010",1449 => X"3C020000",1450 => X"24432278",1451 => X"AC600004",
1452 => X"AC402278",1453 => X"24020011",1454 => X"A0620008",1455 => X"3C023544",
1456 => X"34425441",1457 => X"AF828040",1458 => X"00009825",1459 => X"3C102001",
1460 => X"36103000",1461 => X"3C142001",1462 => X"36943020",1463 => X"24120002",
1464 => X"8F82802C",1465 => X"00000000",1466 => X"14400038",1467 => X"00008825",
1468 => X"AF80802C",1469 => X"A3808030",1470 => X"AF808028",1471 => X"8E020000",
1472 => X"00000000",1473 => X"30420004",1474 => X"10400007",1475 => X"3C032001",
1476 => X"34633000",1477 => X"8C620000",1478 => X"00000000",1479 => X"30420004",
1480 => X"1440FFFC",1481 => X"00000000",1482 => X"8F828040",1483 => X"00000000",
1484 => X"24420001",1485 => X"AF828040",1486 => X"8F848040",1487 => X"0C000544",
1488 => X"00000000",1489 => X"AE820000",1490 => X"AE120000",1491 => X"8E020000",
1492 => X"00000000",1493 => X"30420004",1494 => X"10400007",1495 => X"3C032001",
1496 => X"34633000",1497 => X"8C620000",1498 => X"00000000",1499 => X"30420004",
1500 => X"1440FFFC",1501 => X"00000000",1502 => X"00001825",1503 => X"2402270F",
1504 => X"2442FFFF",1505 => X"0441FFFF",1506 => X"2442FFFF",1507 => X"8F82802C",
1508 => X"00000000",1509 => X"14400005",1510 => X"00000000",1511 => X"24630001",
1512 => X"286203E8",1513 => X"1440FFF6",1514 => X"2402270F",1515 => X"26310001",
1516 => X"2A22000A",1517 => X"10400006",1518 => X"24020001",1519 => X"8F82802C",
1520 => X"00000000",1521 => X"1040FFCA",1522 => X"00000000",1523 => X"24020001",
1524 => X"A3828030",1525 => X"8E020000",1526 => X"00000000",1527 => X"30420004",
1528 => X"10400007",1529 => X"3C032001",1530 => X"34633000",1531 => X"8C620000",
1532 => X"00000000",1533 => X"30420004",1534 => X"1440FFFC",1535 => X"00000000",
1536 => X"0C000581",1537 => X"00000000",1538 => X"AE820000",1539 => X"AE120000",
1540 => X"8E020000",1541 => X"00000000",1542 => X"30420004",1543 => X"10400007",
1544 => X"3C032001",1545 => X"34633000",1546 => X"8C620000",1547 => X"00000000",
1548 => X"30420004",1549 => X"1440FFFC",1550 => X"00000000",1551 => X"00001825",
1552 => X"2402270F",1553 => X"2442FFFF",1554 => X"0441FFFF",1555 => X"2442FFFF",
1556 => X"8F828028",1557 => X"00000000",1558 => X"10400004",1559 => X"00000000",
1560 => X"A3928030",1561 => X"10000009",1562 => X"00000000",1563 => X"24630001",
1564 => X"286203E8",1565 => X"1440FFF3",1566 => X"2402270F",1567 => X"26730001",
1568 => X"2A62000A",1569 => X"1440FF96",1570 => X"00000000",1571 => X"8FBF0024",
1572 => X"8FB40020",1573 => X"8FB3001C",1574 => X"8FB20018",1575 => X"8FB10014",
1576 => X"8FB00010",1577 => X"03E00008",1578 => X"27BD0028",1579 => X"3C022001",
1580 => X"34423000",1581 => X"8C420000",1582 => X"00000000",1583 => X"30420004",
1584 => X"10400008",1585 => X"00000000",1586 => X"3C032001",1587 => X"34633000",
1588 => X"8C620000",1589 => X"00000000",1590 => X"30420004",1591 => X"1440FFFC",
1592 => X"00000000",1593 => X"03E00008",1594 => X"00000000",1595 => X"3C022001",
1596 => X"34423000",1597 => X"8C420000",1598 => X"00000000",1599 => X"30420004",
1600 => X"10400007",1601 => X"3C032001",1602 => X"34633000",1603 => X"8C620000",
1604 => X"00000000",1605 => X"30420004",1606 => X"1440FFFC",1607 => X"00000000",
1608 => X"3C022001",1609 => X"34423020",1610 => X"AC440000",1611 => X"3C032001",
1612 => X"34633000",1613 => X"24020002",1614 => X"03E00008",1615 => X"AC620000",
1616 => X"8F82802C",1617 => X"27BDFFD8",1618 => X"AFBF0020",1619 => X"AFB3001C",
1620 => X"AFB20018",1621 => X"AFB10014",1622 => X"AFB00010",1623 => X"00E09825",
1624 => X"3090FFFF",1625 => X"30B1FFFF",1626 => X"1040003C",1627 => X"30D2FFFF",
1628 => X"0C00062B",1629 => X"00000000",1630 => X"02002025",1631 => X"02202825",
1632 => X"0C0004C4",1633 => X"02403025",1634 => X"3C102001",1635 => X"36103030",
1636 => X"24020806",1637 => X"AE020000",1638 => X"24020001",1639 => X"3C012001",
1640 => X"A4222000",1641 => X"24020800",1642 => X"3C012001",1643 => X"A4222002",
1644 => X"24020604",1645 => X"3C012001",1646 => X"A4222004",1647 => X"24020002",
1648 => X"3C012001",1649 => X"A4222006",1650 => X"3C012001",1651 => X"A4202012",
1652 => X"3C012001",1653 => X"A4202014",1654 => X"3C012001",1655 => X"A4202016",
1656 => X"00131402",1657 => X"3C012001",1658 => X"A4222018",1659 => X"3C012001",
1660 => X"A433201A",1661 => X"3C032001",1662 => X"34630024",1663 => X"8C630000",
1664 => X"3C042001",1665 => X"34840028",1666 => X"8C850000",1667 => X"3C022001",
1668 => X"3442002C",1669 => X"8C420000",1670 => X"3C012001",1671 => X"A422200C",
1672 => X"8F82802C",1673 => X"3C012001",1674 => X"A4232008",1675 => X"8F83802C",
1676 => X"3C012001",1677 => X"A425200A",1678 => X"00021402",1679 => X"3C012001",
1680 => X"A422200E",1681 => X"3C012001",1682 => X"A4232010",1683 => X"0C00063B",
1684 => X"2404002E",1685 => X"24020800",1686 => X"AE020000",1687 => X"8FBF0020",
1688 => X"8FB3001C",1689 => X"8FB20018",1690 => X"8FB10014",1691 => X"8FB00010",
1692 => X"03E00008",1693 => X"27BD0028",1694 => X"27BDFFD8",1695 => X"AFB3001C",
1696 => X"8F938038",1697 => X"24020004",1698 => X"AFBF0020",1699 => X"AFB20018",
1700 => X"AFB10014",1701 => X"AFB00010",1702 => X"AF828038",1703 => X"06600036",
1704 => X"2402FFFF",1705 => X"3C020000",1706 => X"24422340",1707 => X"00131940",
1708 => X"00622021",1709 => X"8C83001C",1710 => X"24020001",1711 => X"14620004",
1712 => X"00000000",1713 => X"3C040000",1714 => X"10000007",1715 => X"24842224",
1716 => X"8C82001C",1717 => X"00000000",1718 => X"14400005",1719 => X"00000000",
1720 => X"3C040000",1721 => X"24842228",1722 => X"0C000099",1723 => X"24050001",
1724 => X"26640030",1725 => X"0C0000D6",1726 => X"308400FF",1727 => X"0C0000D6",
1728 => X"2404000A",1729 => X"3C042001",1730 => X"34843024",1731 => X"8C900000",
1732 => X"3C032001",1733 => X"34633028",1734 => X"8C710000",1735 => X"3C022001",
1736 => X"3442302C",1737 => X"8C520000",1738 => X"3C020000",1739 => X"24422340",
1740 => X"00131940",1741 => X"00621821",1742 => X"8C64000C",1743 => X"8C650010",
1744 => X"8C660014",1745 => X"8C670018",1746 => X"3084FFFF",1747 => X"30A5FFFF",
1748 => X"30C6FFFF",1749 => X"3210FFFF",1750 => X"3231FFFF",1751 => X"0C000650",
1752 => X"3252FFFF",1753 => X"02002025",1754 => X"02202825",1755 => X"0C0004C4",
1756 => X"02403025",1757 => X"2662FFFF",1758 => X"AF828038",1759 => X"8FBF0020",
1760 => X"8FB3001C",1761 => X"8FB20018",1762 => X"8FB10014",1763 => X"8FB00010",
1764 => X"03E00008",1765 => X"27BD0028",1766 => X"27BDFFD0",1767 => X"AFBF002C",
1768 => X"AFB40028",1769 => X"AFB30024",1770 => X"AFB20020",1771 => X"AFB1001C",
1772 => X"AFB00018",1773 => X"2404020A",1774 => X"24053544",1775 => X"0C000490",
1776 => X"24065441",1777 => X"0C0005A2",1778 => X"00000000",1779 => X"3C040000",
1780 => X"2484222C",1781 => X"0C000099",1782 => X"2405000D",1783 => X"8F84802C",
1784 => X"3C100000",1785 => X"26102300",1786 => X"02002825",1787 => X"00009025",
1788 => X"0C00028E",1789 => X"3414EA60",1790 => X"02002025",1791 => X"0C000099",
1792 => X"2405000B",1793 => X"3C040000",1794 => X"2484223C",1795 => X"0C000099",
1796 => X"24050001",1797 => X"3C040000",1798 => X"24842240",1799 => X"0C000099",
1800 => X"24050007",1801 => X"27848028",1802 => X"02002825",1803 => X"0C0001E7",
1804 => X"24060004",1805 => X"02002025",1806 => X"0C000099",1807 => X"24050008",
1808 => X"0C0000D6",1809 => X"2404000A",1810 => X"8F87802C",1811 => X"3404FFFF",
1812 => X"00802825",1813 => X"0C000650",1814 => X"00803025",1815 => X"240470F3",
1816 => X"34059500",1817 => X"0C0004C4",1818 => X"2406721F",1819 => X"3C040000",
1820 => X"0C00026B",1821 => X"24842248",1822 => X"3C030000",1823 => X"24642278",
1824 => X"A0800008",1825 => X"AC602278",1826 => X"8F83802C",1827 => X"00409825",
1828 => X"AC830004",1829 => X"0C00069E",1830 => X"24110400",1831 => X"0C00062B",
1832 => X"3C102001",1833 => X"3610201C",1834 => X"00001825",1835 => X"A2030000",
1836 => X"24630001",1837 => X"0071102A",1838 => X"1440FFFC",1839 => X"26100001",
1840 => X"8F84802C",1841 => X"AFB10010",1842 => X"02602825",1843 => X"00003025",
1844 => X"02543821",1845 => X"30E7FFFF",1846 => X"0C000520",1847 => X"26520001",
1848 => X"0C00063B",1849 => X"00402025",1850 => X"2E420020",1851 => X"1440FFE9",
1852 => X"00000000",1853 => X"0C00069E",1854 => X"00000000",1855 => X"1000FFFD",
1856 => X"00000000",1857 => X"27BDFFA0",1858 => X"AFBF0058",1859 => X"AFB10054",
1860 => X"AFB00050",1861 => X"3C020123",1862 => X"34424567",1863 => X"AC020010",
1864 => X"3C040000",1865 => X"0C000080",1866 => X"24842258",1867 => X"0C0006E6",
1868 => X"00000000",1869 => X"0C00021D",1870 => X"00000000",1871 => X"0C00020A",
1872 => X"00002025",1873 => X"00000000",1874 => X"00000000",1875 => X"00000000",
1876 => X"00000000",1877 => X"00000000",1878 => X"00000000",1879 => X"00000000",
1880 => X"00000000",1881 => X"3C022000",1882 => X"34420070",1883 => X"8C510000",
1884 => X"3C102000",1885 => X"36100060",1886 => X"26310001",1887 => X"AE110000",
1888 => X"00000000",1889 => X"00000000",1890 => X"00000000",1891 => X"00000000",
1892 => X"00000000",1893 => X"00000000",1894 => X"00000000",1895 => X"00000000",
1896 => X"8C510000",1897 => X"3C022000",1898 => X"34420040",1899 => X"AC400000",
1900 => X"3C032000",1901 => X"3463004C",1902 => X"3C020000",1903 => X"24420800",
1904 => X"AC620000",1905 => X"3C032000",1906 => X"34630050",1907 => X"240200FF",
1908 => X"AC620000",1909 => X"0C00001A",1910 => X"24040001",1911 => X"3C040000",
1912 => X"24842268",1913 => X"26310001",1914 => X"0C000080",1915 => X"AE110000",
1916 => X"02202025",1917 => X"27A50010",1918 => X"0C00019B",1919 => X"2406000A",
1920 => X"0C00008E",1921 => X"27A40010",1922 => X"0C0000C4",1923 => X"00000000",
1924 => X"00408825",1925 => X"0C0000D6",1926 => X"322400FF",1927 => X"1000FFFA",
1928 => X"00000000",1929 => X"27BDFFD0",1930 => X"AFBF0028",1931 => X"AFB10024",
1932 => X"AFB00020",1933 => X"00808825",1934 => X"0C00023E",1935 => X"27A50010",
1936 => X"3C040000",1937 => X"24842220",1938 => X"0C000099",1939 => X"24050003",
1940 => X"8FA40010",1941 => X"3C100000",1942 => X"261022C0",1943 => X"2402003B",
1944 => X"A202000B",1945 => X"0C00028E",1946 => X"02002825",1947 => X"02002025",
1948 => X"0C000099",1949 => X"2405000C",1950 => X"8FA40014",1951 => X"0C00028E",
1952 => X"02002825",1953 => X"02002025",1954 => X"0C000099",1955 => X"2405000C",
1956 => X"27A40018",1957 => X"02002825",1958 => X"0C0001E7",1959 => X"24060001",
1960 => X"02002025",1961 => X"0C000099",1962 => X"24050002",1963 => X"0C0000D6",
1964 => X"2404003B",1965 => X"27A40010",1966 => X"3C050000",1967 => X"0C000250",
1968 => X"24A52278",1969 => X"10400019",1970 => X"24020011",1971 => X"93A30018",
1972 => X"00000000",1973 => X"14620006",1974 => X"24020001",1975 => X"02202025",
1976 => X"0C000368",1977 => X"27A50010",1978 => X"10000010",1979 => X"00000000",
1980 => X"14620006",1981 => X"24020006",1982 => X"02202025",1983 => X"0C000326",
1984 => X"27A50010",1985 => X"10000009",1986 => X"00000000",1987 => X"14620005",
1988 => X"02202025",1989 => X"0C000353",1990 => X"27A50010",1991 => X"10000003",
1992 => X"00000000",1993 => X"0C000394",1994 => X"27A50010",1995 => X"8FBF0028",
1996 => X"8FB10024",1997 => X"8FB00020",1998 => X"03E00008",1999 => X"27BD0030",
2000 => X"27BDFFD0",2001 => X"AFBF0028",2002 => X"AFB10024",2003 => X"AFB00020",
2004 => X"3C022001",2005 => X"34425030",2006 => X"00A21026",2007 => X"8C420000",
2008 => X"00808825",2009 => X"3043FFFF",2010 => X"24020800",2011 => X"14620031",
2012 => X"00602025",2013 => X"02202025",2014 => X"0C00023E",2015 => X"27A50010",
2016 => X"3C040000",2017 => X"24842220",2018 => X"0C000099",2019 => X"24050003",
2020 => X"8FA40010",2021 => X"3C100000",2022 => X"261022C0",2023 => X"2402003B",
2024 => X"A202000B",2025 => X"0C00028E",2026 => X"02002825",2027 => X"02002025",
2028 => X"0C000099",2029 => X"2405000C",2030 => X"8FA40014",2031 => X"0C00028E",
2032 => X"02002825",2033 => X"02002025",2034 => X"0C000099",2035 => X"2405000C",
2036 => X"27A40018",2037 => X"02002825",2038 => X"0C0001E7",2039 => X"24060001",
2040 => X"02002025",2041 => X"0C000099",2042 => X"24050002",2043 => X"0C0000D6",
2044 => X"2404003B",2045 => X"27A40010",2046 => X"3C050000",2047 => X"0C000250",
2048 => X"24A52278",2049 => X"1040005B",2050 => X"24020011",2051 => X"93A30018",
2052 => X"00000000",2053 => X"1062003B",2054 => X"24020001",2055 => X"10620040",
2056 => X"24020006",2057 => X"10620045",2058 => X"02202025",2059 => X"10000048",
2060 => X"00000000",2061 => X"24020806",2062 => X"1062004C",2063 => X"2C820600",
2064 => X"1040004C",2065 => X"3C02F000",2066 => X"8E240000",2067 => X"3C034000",
2068 => X"00821024",2069 => X"14430042",2070 => X"3C020001",2071 => X"02202025",
2072 => X"0C00023E",2073 => X"27A50010",2074 => X"3C040000",2075 => X"24842220",
2076 => X"0C000099",2077 => X"24050003",2078 => X"8FA40010",2079 => X"3C100000",
2080 => X"261022C0",2081 => X"2402003B",2082 => X"A202000B",2083 => X"0C00028E",
2084 => X"02002825",2085 => X"02002025",2086 => X"0C000099",2087 => X"2405000C",
2088 => X"8FA40014",2089 => X"0C00028E",2090 => X"02002825",2091 => X"02002025",
2092 => X"0C000099",2093 => X"2405000C",2094 => X"27A40018",2095 => X"02002825",
2096 => X"0C0001E7",2097 => X"24060001",2098 => X"02002025",2099 => X"0C000099",
2100 => X"24050002",2101 => X"0C0000D6",2102 => X"2404003B",2103 => X"27A40010",
2104 => X"3C050000",2105 => X"0C000250",2106 => X"24A52278",2107 => X"10400021",
2108 => X"24020011",2109 => X"93A30018",2110 => X"00000000",2111 => X"14620006",
2112 => X"24020001",2113 => X"02202025",2114 => X"0C000368",2115 => X"27A50010",
2116 => X"10000018",2117 => X"00000000",2118 => X"14620006",2119 => X"24020006",
2120 => X"02202025",2121 => X"0C000326",2122 => X"27A50010",2123 => X"10000011",
2124 => X"00000000",2125 => X"14620006",2126 => X"02202025",2127 => X"02202025",
2128 => X"0C000353",2129 => X"27A50010",2130 => X"1000000A",2131 => X"00000000",
2132 => X"0C000394",2133 => X"27A50010",2134 => X"10000006",2135 => X"00000000",
2136 => X"34420800",2137 => X"14820003",2138 => X"00000000",2139 => X"0C0003AB",
2140 => X"02202025",2141 => X"8FBF0028",2142 => X"8FB10024",2143 => X"8FB00020",
2144 => X"03E00008",2145 => X"27BD0030",2146 => X"00000000",2147 => X"00000000",
2148 => X"00000000",2149 => X"00000000",2150 => X"00000000",2151 => X"00000000",
2152 => X"0A0D0000",2153 => X"5A595857",2154 => X"56555453",2155 => X"5251504F",
2156 => X"4E4D4C4B",2157 => X"4A494847",2158 => X"46454443",2159 => X"42413938",
2160 => X"37363534",2161 => X"33323130",2162 => X"31323334",2163 => X"35363738",
2164 => X"39414243",2165 => X"44454647",2166 => X"48494A4B",2167 => X"4C4D4E4F",
2168 => X"50515253",2169 => X"54555657",2170 => X"58595A00",2171 => X"30313233",
2172 => X"34353637",2173 => X"38394142",2174 => X"43444546",2175 => X"00000000",
2176 => X"0A537461",2177 => X"636B6564",2178 => X"210A0000",2179 => X"443A0000",
2180 => X"433A0000",2181 => X"553A0000",2182 => X"493A0000",2183 => X"0A410000",
2184 => X"0A493A00",2185 => X"61000000",2186 => X"63000000",2187 => X"0A495020",
2188 => X"41646472",2189 => X"6573733A",2190 => X"20000000",2191 => X"3B000000",
2192 => X"4C656173",2193 => X"653A2000",2194 => X"3139322E",2195 => X"3136382E",
2196 => X"3130342E",2197 => X"36340000",2198 => X"48656C6C",2199 => X"6F20576F",
2200 => X"726C640A",2201 => X"00000000",2202 => X"48656C6C",2203 => X"6F20576F",
2204 => X"726C6420",2205 => X"00000000",2206 => X"00000001",2207 => X"00000001",
2208 => X"01000000",2209 => X"2ABCDEF0",2210 => X"20000040",2211 => X"20000044",
2212 => X"2000004C",2213 => X"20000050",2214 => X"00000000",2215 => X"00000000",
2216 => X"00000000",2217 => X"00000000",2218 => X"00000000",2219 => X"FFFFFFFF",
    others => (others => '0')
    );
  signal addr_i : std_logic_vector(M-1 downto 0);

  signal din_i : std_logic_vector(N*8-1 downto 0);

  
begin  -- logic

  din_i <= to_X01(din);


  PROCESS_A : process (clk)
  begin  -- process WRITE_PROCESS
    if rising_edge(clk) then           -- rising clock edge
      addr_i <= addr;
      for i in 0 to N-1 loop
        if wbe(i) = '1' then
          ram(to_integer(unsigned(addr)))(8*i+7 downto 8*i) <= din_i(8*i+7 downto 8*i);
        end if;
      end loop;  -- i
    end if;
  end process PROCESS_A;

  dout <= ram(to_integer(unsigned(addr_i)));

end logic;
