---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_PlasmaBootLoader is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram_PlasmaBootLoader is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"afafafafafafafafaf23ac033c08000cac3c243c241400ac273c243c243c273c",
INIT_01 => X"8f8f8f8f8f8f8f8f8f2300008c8c8c3caf00af00af2340afafafafafafafafaf",
INIT_02 => X"acacacacacacacacacacac40034040033423038f038f8f8f8f8f8f8f8f8f8f8f",
INIT_03 => X"ac303c00100090000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403ac",
INIT_04 => X"02260c9002001a0000afafafaf272703008f240c3c000caf2700030014009024",
INIT_05 => X"8c343c0003001400a024008c001030008d343c353c001827038f8f8f8f020214",
INIT_06 => X"ac033c001430008c343c301030008c343c30038c343c1030008c343c3c143000",
INIT_07 => X"243c353c00243c18ac000001343c01009000243cac03343c24042424ac24343c",
INIT_08 => X"140024ad242404240030002490adad0000912590001400009100243c24353c00",
INIT_09 => X"1800002703008f240c2700a3a300a300af272703008f240c2700a3af27000300",
INIT_0A => X"14002400a0000014303000300000ac8d240424acad2424353c24343c24353c00",
INIT_0B => X"020c02020c323200000000afafafafafaf8faf8faf8faf27ac0324343c000324",
INIT_0C => X"afafaf8f2727038f8f8f8f8f8f8f8f8f000c020c8f021a020c02021a020c021a",
INIT_0D => X"8f000c00240000afaf272703008faf0cafafafaf308f272703008faf0c0030af",
INIT_0E => X"af24afaf272703008f000c000024afaf272703008f000c000024afaf27270300",
INIT_0F => X"000024af24af2727030000000000008f8f93939393270c000024af270c000024",
INIT_10 => X"2727038f8f93000c240c2792240c8e000c92263cafaf27270300008f9393270c",
INIT_11 => X"240c8e000c92263cafaf2727038f8f93000c240c2792240c8e000c92263cafaf",
INIT_12 => X"03008f000c0010243000000c0010243000000caf2727038f8f93000c240c2792",
INIT_13 => X"0000263c000024afafaf93a324a3242414242414002c2c3830a3af0cafaf2727",
INIT_14 => X"240010a32410002c2c3830a3000caf0c278c0000000024afafaf2493af0c008c",
INIT_15 => X"00000090909090ac000000000000909090900003af27038f8f8fa30010a32414",
INIT_16 => X"9090a400009090a400009090a400009090ac00000000000090909090ac000000",
INIT_17 => X"1430932410a71000008f9090a3a3af00000000000027909090909090a4030000",
INIT_18 => X"2424243cafaf18afafafafafafafafaf00272703240010000000973014319324",
INIT_19 => X"00000000af2490242525258f9191912424240024242424242424242424242424",
INIT_1A => X"00000000272726262693929292af000000000000252525252591919191ad0000",
INIT_1B => X"8f8f8f8f8f8f8f8f271400008faf000000000000262626262692929292ae0000",
INIT_1C => X"8f8f8f8f02021402020200028f2400142a020010020000afafafafaf2727038f",
INIT_1D => X"009724142497270c0214020c240002263cafafafafafafafafafaf278f27038f",
INIT_1E => X"0097020c02970200008f00029700240c028f24142c008f24140097241024142c",
INIT_1F => X"00278f2400142a0000008e8e0200100200008e8e000c02278e2626243c020010",
INIT_20 => X"14022626269702140200008e8e001400ac0024028c00243c8e001a0214248e02",
INIT_21 => X"8f27038f8f8f8f8f8f8f8f8f8faf008f000c00000002029700020c02263c8f26",
INIT_22 => X"af8f008f8f020c0000afaf278f002703008f000caf3caf272703008f0000af27",
INIT_23 => X"af2727038f8f8f8f8f00140226ae30a002000c3c001a0000afafafafaf272703",
INIT_24 => X"343c3c1400000c000c243c000c24103cac241030008c343cac24343cac24343c",
INIT_25 => X"000a000000000000001024100024343c00ac2410002400ac343c343c00ac0c24",
INIT_26 => X"00000000000000000000000000000000000000017f00ff0807070e0100000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"a9a8a7a6a5a4a3a2a1bd44e00200000062034202a560a4a0bd1d8404a5059c1c",
INIT_01 => X"a9a8a7a6a5a4a3a2a1a5a086c6c5c406bb00bb00ba5a1abfb9b8afaeadacabaa",
INIT_02 => X"9d9c9e979695949392919084e0029b401bbd60bb60bbbabfb9b8afaeadacabaa",
INIT_03 => X"6242030040008200e000c4e0000085a2e09f9d9c9e979695949392919002e09f",
INIT_04 => X"11100044508020a000b0b1b2bfbdbde000bf8400040000bfbd00e00040008284",
INIT_05 => X"424202c0e00040c543c686e30040420002e707080800a0bde0b0b1b2bf205040",
INIT_06 => X"44e002004042006263038440420042420242e042420240420062630302404200",
INIT_07 => X"42028c0cc24202a062c505406303400042c2420240e042024241420262026303",
INIT_08 => X"40e5e7206363616340424803c22e824800624a488a40e200a2c242020e2909c2",
INIT_09 => X"a00500bde000bf0500a4a0a4a204a204bfbdbde000bf0500a4a0a4bfbd00e000",
INIT_0A => X"40c5c6004382064ac24343420203e002424142eb2c020a08080be7070c290960",
INIT_0B => X"40000060005310e0c0a080b0b1b3b4b5bfb7b7b6b6b2b2bd62e002630300e002",
INIT_0C => X"a7a0bfa2bdbde0b0b1b2b3b4b5b6b7bf00006000a4e0e04000c0a0c040008020",
INIT_0D => X"bf80004004a080a6bfbdbde000bfa200a0a0a0bf84a2bdbde000bfa2000084a0",
INIT_0E => X"b010b0bfbdbde000bfa000a00004a0bfbdbde000bfa000a00004a0bfbdbde000",
INIT_0F => X"a00004a202bfbdbde0454404430302b0bfa5a4a3a2a700a00004b0a700a00004",
INIT_10 => X"bdbde0b0bfa200000500a4060400050000041010b0bfbdbde04302bfa3a2a700",
INIT_11 => X"0400050000041010b0bfbdbde0b0bfa200000500a4060400050000041010b0bf",
INIT_12 => X"e000bf00008062024340000080620283400000bfbdbde0b0bfa200000500a406",
INIT_13 => X"50021010a00004a0a0a082a20282020282020240438342824482b000b1bfbdbd",
INIT_14 => X"0200008202404383428244820000a200a7425002a00004a0a0b11182a200a042",
INIT_15 => X"43030287868382a24746064303028786838200e084bde0b0b1bf910000820282",
INIT_16 => X"8382a362028382a362028382a362028382a247460643030287868382a2474606",
INIT_17 => X"43e2830200a4658202858482a8a7a3666505620203bd888786858283a3e06202",
INIT_18 => X"975e4202a4a5a0b0b1b2b3b4b5b6b7be00bdbde0020200024300838243028302",
INIT_19 => X"43020403a7e7e2c608294aa703244588898a408c8d8e8f589990919253949596",
INIT_1A => X"04430302183910315222032445024544044303026b8cadceef82a3c4e5624544",
INIT_1B => X"b1b2b3b4b5b6b7bede40c700a7c24544044303027394b5d6f782a3c4e5624544",
INIT_1C => X"b1b2b3bf2051403230004060821000400251804032c0a0b0b1b2b3bfbdbde0b0",
INIT_1D => X"00a2026202a3a500004000000540003011b0b1b2b3b4b5b6b7bebfbd82bde0b0",
INIT_1E => X"00a2000055a5a04000820200a240050000a602404200a2026200a30200024042",
INIT_1F => X"40c482100040025243002322c00060436440e483000040c486d4d75602200040",
INIT_20 => X"40a2b5f7d6a2704042430023220040b08382a56563a7e7072200005047072200",
INIT_21 => X"82bde0b0b1b2b3b4b5b6b7bebf8300a3a60006c2024000a2404000001010a694",
INIT_22 => X"82b050bf82000040a0b0bfbd8480bde000bf00008202bfbdbde000bf0040bfbd",
INIT_23 => X"bfbdbde0b0b1b2b3bf00401110424262700000128020a000b0b1b2b3bfbdbde0",
INIT_24 => X"630305e040000000008404000084000462024042004242026202630362026303",
INIT_25 => X"000d000000000000000063408363840400a06340c36300a7c606a50540620002",
INIT_26 => X"00000000000000000000000000000000000000024500ff0406030c0200000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000ff0000200000040020000000ff180015001b0013009300",
INIT_01 => X"00000000000000000000f8200000002000d800d800ff70000000000000000000",
INIT_02 => X"0000000000000000000000600060600000000000000000000000000000000000",
INIT_03 => X"0000200000000000000000002010000000000000000000000000000000000000",
INIT_04 => X"10000000109000888000000000ff00000000120000000000ff000000ff000000",
INIT_05 => X"000020100000ff100000100000000000000020002030000000000000001010ff",
INIT_06 => X"00002000ff0000000020000000000000200000000020ff000000002020000000",
INIT_07 => X"130000206813000000282838002040500010130000000020ffffff0000000020",
INIT_08 => X"ff10000000ffffff400010000000001000000000100010000030130000002058",
INIT_09 => X"0028180000000000000030000012001400ff00000000000000300000ff000000",
INIT_0A => X"ff100018001010000000100010180000ffffff00000000002000002000002030",
INIT_0B => X"28012020000000a888a080000000000000000000000000ff0000000020000000",
INIT_0C => X"00000000ff000000000000000000000000013001002800300028200028012000",
INIT_0D => X"003001280038100000ff000000000001000000000000ff000000000001380000",
INIT_0E => X"00000000ff0000000038013028000000ff0000000038013028000000ff000000",
INIT_0F => X"302800000000ff0000101022101c160000000000000001302800000001302800",
INIT_10 => X"ff000000000000010001000000010000000012000000ff000010120000000001",
INIT_11 => X"00010000000012000000ff000000000000010001000000010000000012000000",
INIT_12 => X"0000000002100000002000021000000020000200ff0000000000000100010000",
INIT_13 => X"101012003028000000008000008000000000000010000000008000020000ff00",
INIT_14 => X"0000008000001000000000800002000100001010302800000000008000013800",
INIT_15 => X"101c160000000000101032101c16000000000000800000000000800000800000",
INIT_16 => X"000000181200000018120000001812000000101032101c160000000000101032",
INIT_17 => X"00008000000000201280000000000018182a18141eff00000000000000001812",
INIT_18 => X"0000150000000000000000000000000030ff000000100010100080ff00008000",
INIT_19 => X"1016221c00000000000000000000000000005800000000000000000000000000",
INIT_1A => X"22101c1600000000000000000000101022101c16000000000000000000001010",
INIT_1B => X"000000000000000000ff10000000101022101c16000000000000000000001010",
INIT_1C => X"000000001080ff108828f82080040000048098001090880000000000ff000000",
INIT_1D => X"00000000000000022000200200f820170000000000000000000000ff80000000",
INIT_1E => X"00002003900028f80080a9200090000320000000200000000000000000000000",
INIT_1F => X"f817800400000480100000008800001818900000980328170000001500f0a800",
INIT_20 => X"ff100000000098ff101000000000ff1000200020001817000028009000000028",
INIT_21 => X"8000000000000000000000000080100030033030302820009028032017000000",
INIT_22 => X"8000100080300128800000ff8010000000000002800000ff0000000000f800ff",
INIT_23 => X"00ff0000000000000000ff100000000018000020980088800000000000ff0000",
INIT_24 => X"0020200038000300021100000411000000000000000000200000002000000020",
INIT_25 => X"000000000000000000ff00ff10008400180000ff100018008400002038000400",
INIT_26 => X"00000000000000000000000000000000000000004c0001020401000400000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"302c2824201c1814109844080012007e4c004c0004fd2a002800400040001301",
INIT_01 => X"302c2824201c181410000924504c400060125c1058fc0054504c4844403c3834",
INIT_02 => X"2824201c1814100c080400000800000801681360115c5854504c4844403c3834",
INIT_03 => X"00ff000009000000080c000810121900082c2824201c1814100c08040000082c",
INIT_04 => X"2a01cf0021250825251014181ce018080010f87900007910e8000800fa000001",
INIT_05 => X"000800250800f52a00012100000808000004000800251120081014181c2521fb",
INIT_06 => X"00080000fc0100000800ff080100000800ff08000400fc080000080000080800",
INIT_07 => X"1c00c400211800280007c025c8002525002114000008c000ffffff010002c000",
INIT_08 => X"e72a010001ffffff25ff04010000000700000100210324000021100001c00021",
INIT_09 => X"21c0252008001803ec1025121103100318e02008001801ec10251018e0000800",
INIT_0A => X"eb2a01250021c30407ff210142400000ffffff00000107c40001c0000fc80025",
INIT_0B => X"25232525e0ffff2525252510141c202430502c48285418c8000802c000000801",
INIT_0C => X"14102038d838081014181c2024282c300063253d4c250425ec252504252e2503",
INIT_0D => X"18259b250325251018e02808002010681c181420ff38d828080020186825ff1c",
INIT_0E => X"10022024d82008001825a92525041018e02008001825a92525061018e0200800",
INIT_0F => X"2525b5100220d8280825210021000020241b1a19181a9b25256510189b252585",
INIT_10 => X"e02008181c100063013d100765230400e007fc00181ce028082500201918189b",
INIT_11 => X"65231000e013fc00181ce02008181c100063013d100b65230800e00bfc00181c",
INIT_12 => X"0800100009250380c025001f250ac0c025000910e82008181c100063013d1013",
INIT_13 => X"2180fc002525061814101320ff1302010280040525010140e011284b2c30c818",
INIT_14 => X"80000813040425010140e011004b1c682000218025256118141001131c682500",
INIT_15 => X"2100001f1e1d1c002121002100001b1a19180008153808282c30130002130204",
INIT_16 => X"31301021002f2e0e21002d2c0c21002b2a082121002100002322212004212100",
INIT_17 => X"0cff1d011006032100191312050400212100210000f805040302010012082100",
INIT_18 => X"130c400000345e080c1014181c20242825d008080380022b26001fff07ff1e02",
INIT_19 => X"21000000002000012020200000000001020325040506070408090a0b08101112",
INIT_1A => X"0021000010202020200000000000212100210000102020202000000000002121",
INIT_1B => X"0c1014181c20242810ba2a003400212100210000102020202000000000002121",
INIT_1C => X"14181c202523f52a21250925150000020123250e2a25251014181c20d8300808",
INIT_1D => X"001e0a76201c10ae257c25e43409254000282c3034383c4044484cb015280810",
INIT_1E => X"001e250e211e2509001540251e25348325140d660000100c6b00200b6f280321",
INIT_1F => X"094015000002012321000c042500282b212500002583254000040c4000252540",
INIT_20 => X"c72a0110101e21db2b21000c0400f52a002104210021400008250d210f010025",
INIT_21 => X"215008282c3034383c4044484c2125102183c021802525222525832540001810",
INIT_22 => X"251021142525b625251014e82525180800100061251810e818080010000910e8",
INIT_23 => X"10e828081014181c2000f72a0100ff002100bd00250c25251014181c20d81808",
INIT_24 => X"600000082500a300ab4800004888050000660508000074000054600000011000",
INIT_25 => X"000000000000000000f101fe2a017f1e250001fe2a0125007f1e600025003fff",
INIT_26 => X"0000000000000000000000000000000000000008460000000000000002000100",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
