-------------------------------------------------------------------------------
-- Inferred BlockRAM with Initial Values
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Ram_PlasmaBootLoader is
  generic (
    N : integer := 4;                -- Width in bytes
    M : integer := 13);               -- Address width

  port (
    clk  : in  std_logic;
    wbe   : in  std_logic_vector(N-1 downto 0)   := (others => '0');
    addr : in  std_logic_vector(M-1 downto 0)   := (others => '0');
    din  : in  std_logic_vector(N*8-1 downto 0) := (others => '0');
    dout : out std_logic_vector(N*8-1 downto 0)
    );

end Ram_PlasmaBootLoader;

architecture logic of Ram_PlasmaBootLoader is

  type mem_file is array(0 to (2**M)-1) of std_logic_vector(N*8-1 downto 0);
  
  signal ram : mem_file := (
    -- Insert initial values below here, eg,
    -- 0 => X"0000",
    -- 1 => X"0001",
    -- <INIT_DATA>
0 => X"3C1C0001",1 => X"279C9343",2 => X"3C050000",3 => X"24A51380",
4 => X"3C040000",5 => X"24841380",6 => X"341D8000",7 => X"ACA00000",
8 => X"00A4182A",9 => X"1460FFFD",10 => X"24A50004",11 => X"3C020000",
12 => X"2442005C",13 => X"3C032000",14 => X"AC62004C",15 => X"0C000489",
16 => X"00000000",17 => X"08000011",18 => X"00000000",19 => X"3C020000",
20 => X"24421380",21 => X"03E00008",22 => X"00000000",23 => X"3C022000",
24 => X"03E00008",25 => X"AC440044",26 => X"40026000",27 => X"03E00008",
28 => X"40846000",29 => X"00000000",30 => X"00000000",31 => X"00000000",
32 => X"23BDFF98",33 => X"AFA10010",34 => X"AFA20014",35 => X"AFA30018",
36 => X"AFA4001C",37 => X"AFA50020",38 => X"AFA60024",39 => X"AFA70028",
40 => X"AFA8002C",41 => X"AFA90030",42 => X"AFAA0034",43 => X"AFAB0038",
44 => X"AFAC003C",45 => X"AFAD0040",46 => X"AFAE0044",47 => X"AFAF0048",
48 => X"AFB8004C",49 => X"AFB90050",50 => X"AFBF0054",51 => X"401A7000",
52 => X"235AFFFC",53 => X"AFBA0058",54 => X"0000D810",55 => X"AFBB005C",
56 => X"0000D812",57 => X"AFBB0060",58 => X"3C062000",59 => X"8CC40040",
60 => X"8CC5004C",61 => X"8CC60050",62 => X"00862024",63 => X"00A0F809",
64 => X"23A50000",65 => X"8FA10010",66 => X"8FA20014",67 => X"8FA30018",
68 => X"8FA4001C",69 => X"8FA50020",70 => X"8FA60024",71 => X"8FA70028",
72 => X"8FA8002C",73 => X"8FA90030",74 => X"8FAA0034",75 => X"8FAB0038",
76 => X"8FAC003C",77 => X"8FAD0040",78 => X"8FAE0044",79 => X"8FAF0048",
80 => X"8FB8004C",81 => X"8FB90050",82 => X"8FBF0054",83 => X"8FBA0058",
84 => X"8FBB005C",85 => X"03600011",86 => X"8FBB0060",87 => X"03600013",
88 => X"23BD0068",89 => X"341B0001",90 => X"03400008",91 => X"409B6000",
92 => X"AC900000",93 => X"AC910004",94 => X"AC920008",95 => X"AC93000C",
96 => X"AC940010",97 => X"AC950014",98 => X"AC960018",99 => X"AC97001C",
100 => X"AC9E0020",101 => X"AC9C0024",102 => X"AC9D0028",103 => X"AC9F002C",
104 => X"03E00008",105 => X"34020000",106 => X"8C900000",107 => X"8C910004",
108 => X"8C920008",109 => X"8C93000C",110 => X"8C940010",111 => X"8C950014",
112 => X"8C960018",113 => X"8C97001C",114 => X"8C9E0020",115 => X"8C9C0024",
116 => X"8C9D0028",117 => X"8C9F002C",118 => X"03E00008",119 => X"34A20000",
120 => X"00850019",121 => X"00001012",122 => X"00002010",123 => X"03E00008",
124 => X"ACC40000",125 => X"0000000C",126 => X"03E00008",127 => X"00000000",
128 => X"90820000",129 => X"00000000",130 => X"10400009",131 => X"00000000",
132 => X"3C032000",133 => X"304200FF",134 => X"AC620000",135 => X"24840001",
136 => X"90820000",137 => X"00000000",138 => X"1440FFFA",139 => X"00000000",
140 => X"03E00008",141 => X"00000000",142 => X"27BDFFE8",143 => X"AFBF0010",
144 => X"0C000080",145 => X"00000000",146 => X"3C040000",147 => X"0C000080",
148 => X"24841328",149 => X"8FBF0010",150 => X"00000000",151 => X"03E00008",
152 => X"27BD0018",153 => X"27BDFFE0",154 => X"AFBF001C",155 => X"AFB20018",
156 => X"AFB10014",157 => X"AFB00010",158 => X"00008025",159 => X"00A08825",
160 => X"1A200008",161 => X"00809025",162 => X"02501021",163 => X"90440000",
164 => X"0C0000D6",165 => X"26100001",166 => X"0211102A",167 => X"1440FFFB",
168 => X"02501021",169 => X"02201025",170 => X"8FBF001C",171 => X"8FB20018",
172 => X"8FB10014",173 => X"8FB00010",174 => X"03E00008",175 => X"27BD0020",
176 => X"18A00011",177 => X"00003025",178 => X"3C082000",179 => X"35080008",
180 => X"3C072000",181 => X"34E70004",182 => X"8D020000",183 => X"00000000",
184 => X"30420008",185 => X"10400008",186 => X"00000000",187 => X"8CE30000",
188 => X"00861021",189 => X"24C60001",190 => X"A0430000",191 => X"00C5102A",
192 => X"1440FFF5",193 => X"00000000",194 => X"03E00008",195 => X"00C01025",
196 => X"3C022000",197 => X"34420008",198 => X"8C420000",199 => X"00000000",
200 => X"30420008",201 => X"14400008",202 => X"3C022000",203 => X"3C032000",
204 => X"34630008",205 => X"8C620000",206 => X"00000000",207 => X"30420008",
208 => X"1040FFFC",209 => X"3C022000",210 => X"34420004",211 => X"8C420000",
212 => X"03E00008",213 => X"304200FF",214 => X"3C022000",215 => X"34420008",
216 => X"8C420000",217 => X"00000000",218 => X"30420001",219 => X"10400008",
220 => X"308400FF",221 => X"3C032000",222 => X"34630008",223 => X"8C620000",
224 => X"00000000",225 => X"30420001",226 => X"1440FFFC",227 => X"00000000",
228 => X"3C022000",229 => X"03E00008",230 => X"AC440000",231 => X"3C032000",
232 => X"346300C0",233 => X"24020002",234 => X"AC620000",235 => X"24020001",
236 => X"2442FFFF",237 => X"0441FFFF",238 => X"2442FFFF",239 => X"3C022000",
240 => X"344200C0",241 => X"03E00008",242 => X"AC400000",243 => X"3C020000",
244 => X"24421344",245 => X"00C21021",246 => X"90420000",247 => X"00005025",
248 => X"01404025",249 => X"3C032000",250 => X"346300C8",251 => X"01403825",
252 => X"000528C0",253 => X"00C52807",254 => X"AC620000",255 => X"18A00028",
256 => X"3C020000",257 => X"24421348",258 => X"00C26821",259 => X"3C0C2000",
260 => X"358C00C4",261 => X"3C020000",262 => X"2442134C",263 => X"00C25821",
264 => X"3C092000",265 => X"352900C0",266 => X"240E0001",267 => X"3C020000",
268 => X"24421340",269 => X"00C23021",270 => X"91A20000",271 => X"00000000",
272 => X"00E21024",273 => X"14400003",274 => X"008A1021",275 => X"90480000",
276 => X"254A0001",277 => X"91620000",278 => X"00000000",279 => X"00481007",
280 => X"AD820000",281 => X"AD2E0000",282 => X"90C20000",283 => X"24030001",
284 => X"00481004",285 => X"304200FF",286 => X"00404025",287 => X"2463FFFF",
288 => X"0461FFFF",289 => X"2463FFFF",290 => X"24630001",291 => X"AD200000",
292 => X"24E70001",293 => X"00E5102A",294 => X"1440FFE7",295 => X"00000000",
296 => X"03E00008",297 => X"00000000",298 => X"27BDFFE0",299 => X"AFBF0018",
300 => X"A3A40010",301 => X"00A03025",302 => X"27A40010",303 => X"0C0000F3",
304 => X"24050001",305 => X"8FBF0018",306 => X"00000000",307 => X"03E00008",
308 => X"27BD0020",309 => X"27BDFFE0",310 => X"AFBF0018",311 => X"00041403",
312 => X"A3A20010",313 => X"00041203",314 => X"A3A20011",315 => X"A3A40012",
316 => X"00A03025",317 => X"27A40010",318 => X"0C0000F3",319 => X"24050003",
320 => X"8FBF0018",321 => X"00000000",322 => X"03E00008",323 => X"27BD0020",
324 => X"00001825",325 => X"000528C0",326 => X"18A00021",327 => X"00603025",
328 => X"3C092000",329 => X"352900C8",330 => X"240C000F",331 => X"3C072000",
332 => X"34E700C0",333 => X"240B0001",334 => X"3C082000",335 => X"350800C4",
336 => X"240A0007",337 => X"24020001",338 => X"AD2C0000",339 => X"ACEB0000",
340 => X"2442FFFF",341 => X"0441FFFF",342 => X"2442FFFF",343 => X"8D020000",
344 => X"ACE00000",345 => X"00031840",346 => X"00021042",347 => X"30420001",
348 => X"00431021",349 => X"304300FF",350 => X"30C20007",351 => X"144A0004",
352 => X"000610C3",353 => X"00821021",354 => X"A0430000",355 => X"00001825",
356 => X"24C60001",357 => X"00C5102A",358 => X"1440FFEB",359 => X"24020001",
360 => X"03E00008",361 => X"00000000",362 => X"3C032000",363 => X"346300C0",
364 => X"24020002",365 => X"03E00008",366 => X"AC620000",367 => X"27BDFFC8",
368 => X"AFB20018",369 => X"8FB20054",370 => X"AFB60028",371 => X"8FB60048",
372 => X"AFB7002C",373 => X"8FB70050",374 => X"AFBF0030",375 => X"AFB50024",
376 => X"AFB40020",377 => X"AFB3001C",378 => X"AFB10014",379 => X"AFB00010",
380 => X"00808025",381 => X"00A0A025",382 => X"00C08825",383 => X"00E0A825",
384 => X"321000FF",385 => X"325300FF",386 => X"0C0000E7",387 => X"02602025",
388 => X"02002025",389 => X"0C00012A",390 => X"02402825",391 => X"1A200003",
392 => X"02802025",393 => X"0C000135",394 => X"02402825",395 => X"1AC00004",
396 => X"02A02025",397 => X"02C02825",398 => X"0C0000F3",399 => X"02403025",
400 => X"1AE00004",401 => X"02E02825",402 => X"8FA4004C",403 => X"0C000144",
404 => X"02603025",405 => X"0C00016A",406 => X"00000000",407 => X"8FBF0030",
408 => X"8FB7002C",409 => X"8FB60028",410 => X"8FB50024",411 => X"8FB40020",
412 => X"8FB3001C",413 => X"8FB20018",414 => X"8FB10014",415 => X"8FB00010",
416 => X"03E00008",417 => X"27BD0038",418 => X"27BDFFD8",419 => X"8FA20038",
420 => X"AFBF0020",421 => X"AFA00010",422 => X"AFA70014",423 => X"AFA0001C",
424 => X"308400FF",425 => X"00003825",426 => X"0C00016F",427 => X"AFA20018",
428 => X"8FBF0020",429 => X"00000000",430 => X"03E00008",431 => X"27BD0028",
432 => X"27BDFFD8",433 => X"8FA20038",434 => X"308400FF",435 => X"AFBF0020",
436 => X"AFA00014",437 => X"AFA00018",438 => X"AFA0001C",439 => X"0C00016F",
440 => X"AFA20010",441 => X"8FBF0020",442 => X"00000000",443 => X"03E00008",
444 => X"27BD0028",445 => X"27BDFFE0",446 => X"AFBF0018",447 => X"AFA60010",
448 => X"00801025",449 => X"00A03825",450 => X"24040003",451 => X"00402825",
452 => X"0C0001A2",453 => X"00803025",454 => X"8FBF0018",455 => X"00000000",
456 => X"03E00008",457 => X"27BD0020",458 => X"27BDFFE0",459 => X"AFBF0018",
460 => X"AFA00010",461 => X"24040006",462 => X"00002825",463 => X"00A03025",
464 => X"0C0001B0",465 => X"00A03825",466 => X"8FBF0018",467 => X"00000000",
468 => X"03E00008",469 => X"27BD0020",470 => X"27BDFFE0",471 => X"AFBF0018",
472 => X"AFA00010",473 => X"24040004",474 => X"00002825",475 => X"00A03025",
476 => X"0C0001B0",477 => X"00A03825",478 => X"8FBF0018",479 => X"00000000",
480 => X"03E00008",481 => X"27BD0020",482 => X"27BDFFD8",483 => X"AFBF0024",
484 => X"AFB00020",485 => X"24100002",486 => X"AFB00010",487 => X"24040085",
488 => X"00002825",489 => X"00A03025",490 => X"0C0001A2",491 => X"27A70018",
492 => X"AFB00010",493 => X"24040065",494 => X"00002825",495 => X"00A03025",
496 => X"0C0001A2",497 => X"27A7001A",498 => X"93A20018",499 => X"93A30019",
500 => X"93A4001A",501 => X"93A5001B",502 => X"8FBF0024",503 => X"8FB00020",
504 => X"00021600",505 => X"00031C00",506 => X"00431021",507 => X"00042200",
508 => X"00441021",509 => X"00451025",510 => X"03E00008",511 => X"27BD0028",
512 => X"27BDFFD8",513 => X"AFBF0020",514 => X"24020002",515 => X"AFA20010",
516 => X"240400B5",517 => X"00002825",518 => X"00A03025",519 => X"0C0001A2",
520 => X"27A70018",521 => X"93A20018",522 => X"93A30019",523 => X"8FBF0020",
524 => X"00021200",525 => X"00431025",526 => X"03E00008",527 => X"27BD0028",
528 => X"27BDFFE0",529 => X"AFBF001C",530 => X"AFB00018",531 => X"3C100000",
532 => X"2610132C",533 => X"92040007",534 => X"0C0000E7",535 => X"00000000",
536 => X"8E050004",537 => X"0C00012A",538 => X"24040065",539 => X"92060007",
540 => X"27A40010",541 => X"0C000144",542 => X"24050001",543 => X"0C00016A",
544 => X"00000000",545 => X"93A20010",546 => X"8FBF001C",547 => X"8FB00018",
548 => X"03E00008",549 => X"27BD0020",550 => X"27BDFFE0",551 => X"AFBF001C",
552 => X"AFB00018",553 => X"3C100000",554 => X"2610132C",555 => X"9204000B",
556 => X"0C0000E7",557 => X"00000000",558 => X"8E050008",559 => X"0C00012A",
560 => X"24040065",561 => X"9206000B",562 => X"27A40010",563 => X"0C000144",
564 => X"24050001",565 => X"0C00016A",566 => X"00000000",567 => X"93A20010",
568 => X"8FBF001C",569 => X"8FB00018",570 => X"03E00008",571 => X"27BD0020",
572 => X"27BDFFE0",573 => X"AFBF001C",574 => X"AFB00018",575 => X"3C100000",
576 => X"2610132C",577 => X"92040013",578 => X"0C0000E7",579 => X"00000000",
580 => X"8E050010",581 => X"0C00012A",582 => X"24040065",583 => X"92060013",
584 => X"27A40010",585 => X"0C000144",586 => X"24050001",587 => X"0C00016A",
588 => X"00000000",589 => X"93A20010",590 => X"8FBF001C",591 => X"8FB00018",
592 => X"03E00008",593 => X"27BD0020",594 => X"27BDFFE8",595 => X"AFBF0010",
596 => X"0C000210",597 => X"00000000",598 => X"00402025",599 => X"308300C0",
600 => X"240200C0",601 => X"1062000A",602 => X"00801025",603 => X"0C000226",
604 => X"00000000",605 => X"00402025",606 => X"304300C0",607 => X"24020080",
608 => X"10620003",609 => X"00801025",610 => X"0C000210",611 => X"00000000",
612 => X"8FBF0010",613 => X"00000000",614 => X"03E00008",615 => X"27BD0018",
616 => X"27BDFFC8",617 => X"AFBF0030",618 => X"AFB1002C",619 => X"0C000252",
620 => X"AFB00028",621 => X"A3828025",622 => X"304400E0",623 => X"38820040",
624 => X"2C420001",625 => X"2C830001",626 => X"00431025",627 => X"14400005",
628 => X"24020004",629 => X"24020080",630 => X"14820002",631 => X"24020001",
632 => X"24020002",633 => X"A3828027",634 => X"240200FF",635 => X"A3A20020",
636 => X"93828027",637 => X"AFA00010",638 => X"AFA00014",639 => X"AFA00018",
640 => X"24040006",641 => X"00002825",642 => X"00A03025",643 => X"3C100000",
644 => X"2610132C",645 => X"00021080",646 => X"00501021",647 => X"8C420000",
648 => X"00A03825",649 => X"0C00016F",650 => X"AFA2001C",651 => X"93828027",
652 => X"24110001",653 => X"AFB10010",654 => X"AFA00014",655 => X"AFA00018",
656 => X"24040061",657 => X"00002825",658 => X"00A03025",659 => X"00021080",
660 => X"00501021",661 => X"8C420000",662 => X"27A70020",663 => X"0C00016F",
664 => X"AFA2001C",665 => X"0C000252",666 => X"00000000",667 => X"A3828025",
668 => X"304400E0",669 => X"38820040",670 => X"2C420001",671 => X"2C830001",
672 => X"00431025",673 => X"10400004",674 => X"24020004",675 => X"A3828027",
676 => X"10000008",677 => X"00000000",678 => X"24020080",679 => X"14820004",
680 => X"24020002",681 => X"A3828027",682 => X"10000002",683 => X"00000000",
684 => X"A3918027",685 => X"8FBF0030",686 => X"8FB1002C",687 => X"8FB00028",
688 => X"03E00008",689 => X"27BD0038",690 => X"AF848029",691 => X"03E00008",
692 => X"00000000",693 => X"90820018",694 => X"90830019",695 => X"9086001A",
696 => X"9087001B",697 => X"00021600",698 => X"00031C00",699 => X"00431021",
700 => X"00063200",701 => X"00461021",702 => X"00471021",703 => X"ACA20000",
704 => X"9082001C",705 => X"9083001D",706 => X"9086001E",707 => X"9087001F",
708 => X"00021600",709 => X"00031C00",710 => X"00431021",711 => X"00063200",
712 => X"00461021",713 => X"00471021",714 => X"ACA20004",715 => X"90820020",
716 => X"90830021",717 => X"90860022",718 => X"90870023",719 => X"00021600",
720 => X"00031C00",721 => X"00431021",722 => X"00063200",723 => X"00461021",
724 => X"00471021",725 => X"ACA20008",726 => X"9082002A",727 => X"9083002B",
728 => X"00021200",729 => X"00621821",730 => X"A4A3000C",731 => X"9082002C",
732 => X"9083002D",733 => X"00021200",734 => X"00621821",735 => X"A4A3000E",
736 => X"9082002E",737 => X"9083002F",738 => X"00021200",739 => X"00621821",
740 => X"A4A30010",741 => X"90820030",742 => X"90830031",743 => X"00021200",
744 => X"00621821",745 => X"03E00008",746 => X"A4A30012",747 => X"90830000",
748 => X"90820001",749 => X"90850002",750 => X"90860003",751 => X"90870004",
752 => X"90880005",753 => X"27BDFFF8",754 => X"00031E00",755 => X"00021400",
756 => X"00621821",757 => X"00052A00",758 => X"00651821",759 => X"00661821",
760 => X"AFA30000",761 => X"A3A70004",762 => X"A3A80005",763 => X"90820012",
764 => X"90840013",765 => X"8F85802D",766 => X"00021200",767 => X"00822021",
768 => X"10650003",769 => X"A7A40006",770 => X"10000010",771 => X"24020001",
772 => X"93838031",773 => X"30E200FF",774 => X"1443000C",775 => X"24020002",
776 => X"93838032",777 => X"310200FF",778 => X"14430007",779 => X"3082FFFF",
780 => X"97838033",781 => X"00000000",782 => X"00431026",783 => X"0002102B",
784 => X"10000002",785 => X"00021080",786 => X"24020003",787 => X"03E00008",
788 => X"27BD0008",789 => X"27BDFFD0",790 => X"00003825",791 => X"AFBE0028",
792 => X"AFB70024",793 => X"AFB60020",794 => X"AFB5001C",795 => X"AFB40018",
796 => X"AFB30014",797 => X"AFB20010",798 => X"AFB1000C",799 => X"AFB00008",
800 => X"18A0005B",801 => X"AFA50034",802 => X"AFA40000",803 => X"24DE000C",
804 => X"24970013",805 => X"24960012",806 => X"24950011",807 => X"24940010",
808 => X"24D30008",809 => X"2492000B",810 => X"2491000A",811 => X"24900009",
812 => X"24990008",813 => X"24D80004",814 => X"248F0007",815 => X"248E0006",
816 => X"248D0005",817 => X"248C0004",818 => X"248B0003",819 => X"248A0002",
820 => X"24890001",821 => X"91650000",822 => X"91440000",823 => X"91230000",
824 => X"8FA80000",825 => X"256B0020",826 => X"254A0020",827 => X"25290020",
828 => X"24E70001",829 => X"91020000",830 => X"25080020",831 => X"AFA80000",
832 => X"00031C00",833 => X"00042200",834 => X"00021600",835 => X"00431021",
836 => X"00441021",837 => X"00451021",838 => X"ACC20000",839 => X"91E50000",
840 => X"91C40000",841 => X"91A30000",842 => X"91820000",843 => X"25EF0020",
844 => X"25CE0020",845 => X"25AD0020",846 => X"258C0020",847 => X"24C60010",
848 => X"00021600",849 => X"00031C00",850 => X"00431021",851 => X"00042200",
852 => X"00441021",853 => X"00451021",854 => X"AF020000",855 => X"92450000",
856 => X"92240000",857 => X"92030000",858 => X"93220000",859 => X"26520020",
860 => X"26310020",861 => X"26100020",862 => X"27390020",863 => X"27180010",
864 => X"00021600",865 => X"00031C00",866 => X"00431021",867 => X"00042200",
868 => X"00441021",869 => X"00451021",870 => X"AE620000",871 => X"92E50000",
872 => X"92C40000",873 => X"92A30000",874 => X"92820000",875 => X"26F70020",
876 => X"26D60020",877 => X"26B50020",878 => X"26940020",879 => X"26730010",
880 => X"00021600",881 => X"00031C00",882 => X"00431021",883 => X"00042200",
884 => X"00441021",885 => X"00451021",886 => X"AFC20000",887 => X"8FA80034",
888 => X"00000000",889 => X"00E8102A",890 => X"1440FFBA",891 => X"27DE0010",
892 => X"8FBE0028",893 => X"8FB70024",894 => X"8FB60020",895 => X"8FB5001C",
896 => X"8FB40018",897 => X"8FB30014",898 => X"8FB20010",899 => X"8FB1000C",
900 => X"8FB00008",901 => X"03E00008",902 => X"27BD0030",903 => X"27BDFFD8",
904 => X"AFBF0020",905 => X"AFB3001C",906 => X"AFB20018",907 => X"AFB10014",
908 => X"AFB00010",909 => X"00A08825",910 => X"00C09025",911 => X"0232102A",
912 => X"1040000E",913 => X"00809825",914 => X"02518023",915 => X"2A020401",
916 => X"14400002",917 => X"00000000",918 => X"24100400",919 => X"8F828029",
920 => X"02602025",921 => X"0040F809",922 => X"02002825",923 => X"02308821",
924 => X"0232102A",925 => X"1440FFF5",926 => X"02518023",927 => X"02201025",
928 => X"8FBF0020",929 => X"8FB3001C",930 => X"8FB20018",931 => X"8FB10014",
932 => X"8FB00010",933 => X"03E00008",934 => X"27BD0028",935 => X"8F828029",
936 => X"27BDF9A8",937 => X"AFBF0654",938 => X"AFBE0650",939 => X"AFB7064C",
940 => X"AFB60648",941 => X"AFB50644",942 => X"AFB40640",943 => X"AFB3063C",
944 => X"AFB20638",945 => X"AFB10634",946 => X"AFB00630",947 => X"27B00028",
948 => X"02002025",949 => X"0040F809",950 => X"24050034",951 => X"0C0002EB",
952 => X"02002025",953 => X"1440007F",954 => X"02002025",955 => X"0C0002B5",
956 => X"27A50010",957 => X"97A3001C",958 => X"24020020",959 => X"14620079",
960 => X"24020005",961 => X"97A2001E",962 => X"00000000",963 => X"2C420021",
964 => X"14400003",965 => X"24020028",966 => X"10000072",967 => X"24020006",
968 => X"97A30020",969 => X"00000000",970 => X"10620005",971 => X"24020007",
972 => X"1000006C",973 => X"00000000",974 => X"1000006A",975 => X"24020008",
976 => X"8FA60014",977 => X"02002025",978 => X"0C000387",979 => X"24050034",
980 => X"00409025",981 => X"97A2001E",982 => X"02002025",983 => X"0002A140",
984 => X"8F828029",985 => X"00000000",986 => X"0040F809",987 => X"02802825",
988 => X"97A5001E",989 => X"02549021",990 => X"02002025",991 => X"27B10428",
992 => X"0C000315",993 => X"02203025",994 => X"97A2001E",995 => X"00000000",
996 => X"10400043",997 => X"0000A025",998 => X"AFB00628",999 => X"0220F025",
1000 => X"27B70434",1001 => X"27B5042C",1002 => X"27B60430",1003 => X"8EC20000",
1004 => X"00000000",1005 => X"2C422000",1006 => X"1440FFDF",1007 => X"27A40028",
1008 => X"8EA60000",1009 => X"02402825",1010 => X"0C000387",1011 => X"00009825",
1012 => X"8EA30000",1013 => X"8EE40000",1014 => X"00409025",1015 => X"00641821",
1016 => X"0243182B",1017 => X"10600026",1018 => X"00000000",1019 => X"03C08825",
1020 => X"8E220004",1021 => X"8E23000C",1022 => X"00000000",1023 => X"00431021",
1024 => X"00528023",1025 => X"2A020401",1026 => X"14400002",1027 => X"00000000",
1028 => X"24100400",1029 => X"8F828029",1030 => X"27A40028",1031 => X"0040F809",
1032 => X"02002825",1033 => X"8E220000",1034 => X"24070001",1035 => X"1447000D",
1036 => X"02509021",1037 => X"1A00000B",1038 => X"00002825",1039 => X"8FA70628",
1040 => X"8E220008",1041 => X"02652021",1042 => X"00E51821",1043 => X"90630000",
1044 => X"24A50001",1045 => X"00822021",1046 => X"00B0102A",1047 => X"1440FFF7",
1048 => X"A0830000",1049 => X"8E220004",1050 => X"8E23000C",1051 => X"00000000",
1052 => X"00431021",1053 => X"0242102B",1054 => X"1440FFDD",1055 => X"02709821",
1056 => X"97A2001E",1057 => X"27DE0010",1058 => X"26F70010",1059 => X"26B50010",
1060 => X"26940001",1061 => X"0282102A",1062 => X"1440FFC4",1063 => X"26D60010",
1064 => X"8FA60018",1065 => X"27B00028",1066 => X"02002025",1067 => X"0C000387",
1068 => X"02402825",1069 => X"00409025",1070 => X"97A20022",1071 => X"02002025",
1072 => X"02402825",1073 => X"00023080",1074 => X"00C23021",1075 => X"000630C0",
1076 => X"0C000387",1077 => X"00A63021",1078 => X"8FA30010",1079 => X"00001025",
1080 => X"AF838035",1081 => X"8FBF0654",1082 => X"8FBE0650",1083 => X"8FB7064C",
1084 => X"8FB60648",1085 => X"8FB50644",1086 => X"8FB40640",1087 => X"8FB3063C",
1088 => X"8FB20638",1089 => X"8FB10634",1090 => X"8FB00630",1091 => X"03E00008",
1092 => X"27BD0658",1093 => X"8F828035",1094 => X"27BDFFE8",1095 => X"AFBF0010",
1096 => X"0040F809",1097 => X"00000000",1098 => X"8FBF0010",1099 => X"00000000",
1100 => X"03E00008",1101 => X"27BD0018",1102 => X"27BDFFE8",1103 => X"AFBF0010",
1104 => X"3C020018",1105 => X"AF828039",1106 => X"0C000268",1107 => X"00000000",
1108 => X"8FBF0010",1109 => X"00000000",1110 => X"03E00008",1111 => X"27BD0018",
1112 => X"3C032000",1113 => X"34630010",1114 => X"24020001",1115 => X"03E00008",
1116 => X"AC620000",1117 => X"00801025",1118 => X"8F848039",1119 => X"27BDFFE8",
1120 => X"AFBF0014",1121 => X"AFB00010",1122 => X"00A08025",1123 => X"00402825",
1124 => X"0C0001BD",1125 => X"02003025",1126 => X"8F828039",1127 => X"8FBF0014",
1128 => X"00501021",1129 => X"8FB00010",1130 => X"AF828039",1131 => X"03E00008",
1132 => X"27BD0018",1133 => X"27BDFFD8",1134 => X"AFBF0020",1135 => X"AFB3001C",
1136 => X"AFB20018",1137 => X"AFB10014",1138 => X"AFB00010",1139 => X"00008025",
1140 => X"00A08825",1141 => X"1A20000C",1142 => X"00809825",1143 => X"3C122000",
1144 => X"0C0000C4",1145 => X"00000000",1146 => X"02701821",1147 => X"A0620000",
1148 => X"304200FF",1149 => X"AE420000",1150 => X"26100001",1151 => X"0211102A",
1152 => X"1440FFF7",1153 => X"00000000",1154 => X"8FBF0020",1155 => X"8FB3001C",
1156 => X"8FB20018",1157 => X"8FB10014",1158 => X"8FB00010",1159 => X"03E00008",
1160 => X"27BD0028",1161 => X"27BDFFE8",1162 => X"AFBF0010",1163 => X"3C022000",
1164 => X"34420074",1165 => X"8C420000",1166 => X"00000000",1167 => X"30420008",
1168 => X"10400008",1169 => X"3C022000",1170 => X"34420060",1171 => X"24030066",
1172 => X"0C000458",1173 => X"AC430000",1174 => X"3C040000",1175 => X"10000007",
1176 => X"248411B4",1177 => X"34420060",1178 => X"24030054",1179 => X"0C00044E",
1180 => X"AC430000",1181 => X"3C040000",1182 => X"24841174",1183 => X"0C0002B2",
1184 => X"00000000",1185 => X"0C0003A7",1186 => X"00000000",1187 => X"00403825",
1188 => X"14E0000C",1189 => X"3C052000",1190 => X"3C032000",1191 => X"34630060",
1192 => X"240200FF",1193 => X"0C000013",1194 => X"AC620000",1195 => X"8F838011",
1196 => X"2442FFFF",1197 => X"0C000445",1198 => X"AC620000",1199 => X"00403825",
1200 => X"3C052000",1201 => X"34A50060",1202 => X"3C06001E",1203 => X"34C6847F",
1204 => X"ACA70000",1205 => X"00001825",1206 => X"24630001",1207 => X"00C3102A",
1208 => X"1040FFFE",1209 => X"24630001",1210 => X"ACA00000",1211 => X"00001825",
1212 => X"3C04001E",1213 => X"3484847F",1214 => X"24630001",1215 => X"0083102A",
1216 => X"1040FFFE",1217 => X"24630001",1218 => X"1000FFF1",1219 => X"00000000",
1220 => X"00000000",1221 => X"00000000",1222 => X"00000000",1223 => X"00000000",
1224 => X"00000000",1225 => X"00000000",1226 => X"0A0D0000",1227 => X"00000000",
1228 => X"00000000",1229 => X"00000001",1230 => X"00000000",1231 => X"00000002",
1232 => X"01020400",1233 => X"0E0C0000",1234 => X"07030100",1235 => X"07060400",
1236 => X"08040200",1237 => X"2ABCDEF0",1238 => X"20000040",1239 => X"20000044",
1240 => X"2000004C",1241 => X"20000050",1242 => X"FFFF0100",1243 => X"00000000",
1244 => X"7F454C46",1245 => X"01020008",1246 => X"00000000",1247 => X"00000000",
    others => (others => '0')
    );
  signal addr_i : std_logic_vector(M-1 downto 0);

  signal din_i : std_logic_vector(N*8-1 downto 0);

  
begin  -- logic

  din_i <= to_X01(din);


  PROCESS_A : process (clk)
  begin  -- process WRITE_PROCESS
    if rising_edge(clk) then           -- rising clock edge
      addr_i <= addr;
      for i in 0 to N-1 loop
        if wbe(i) = '1' then
          ram(to_integer(unsigned(addr)))(8*i+7 downto 8*i) <= din_i(8*i+7 downto 8*i);
        end if;
      end loop;  -- i
    end if;
  end process PROCESS_A;

  dout <= ram(to_integer(unsigned(addr_i)));

end logic;
