---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_PlasmaBootLoader is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram_PlasmaBootLoader is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"000000400340ac033c0003243c0008000cac3c243c241400ac34243c243c273c",
INIT_01 => X"00008c8c8c3caf00af00af2340afafafafafafafafafafafafafafafafafaf23",
INIT_02 => X"acacacac40033423038f038f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f23",
INIT_03 => X"000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403acacacacacacacac",
INIT_04 => X"0000afafafaf272703008f240c3c000caf2700030014009024ac303c00100090",
INIT_05 => X"00a024008c001030008d343c353c001827038f8f8f8f02021402260c9002001a",
INIT_06 => X"8c343c301030008c343c30038c343c1030008c343c3c1430008c343c00030014",
INIT_07 => X"18ac000001343c01009000243cac03343c24042424ac24343cac033c00143000",
INIT_08 => X"240030002490adad0000912590001400009100243c24353c00243c353c00243c",
INIT_09 => X"240c2700a3a300a300af272703008f240c2700a3af27000300140024ad242404",
INIT_0A => X"14303000300000ac8d240424acad2424353c24343c24353c001800002703008f",
INIT_0B => X"00000000afafafafafaf8faf8faf8faf27ac0324343c00032414002400a00000",
INIT_0C => X"8f8f8f8f8f8f8f8f8f000c020c8f021a020c02021a020c021a020c02020c3232",
INIT_0D => X"afaf272703008faf0cafafafaf308f272703008faf0c0030afafafaf8f272703",
INIT_0E => X"008f000c000024afaf272703008f000c000024afaf272703008f000c00240000",
INIT_0F => X"27030000000000008f8f93939393270c000024af270c000024af24afaf272703",
INIT_10 => X"0c240c2792240c8e000c92263cafaf27270300008f9393270c000024af24af27",
INIT_11 => X"3cafaf2727038f8f93000c240c2792240c8e000c92263cafaf2727038f8f9300",
INIT_12 => X"243000000c0010243000000caf2727038f8f93000c240c2792240c8e000c9226",
INIT_13 => X"afafaf93a324a3242414242414002c2c3830a3af0cafaf272703008f000c0010",
INIT_14 => X"2c2c3830a3000caf0c278c0000000024afafaf2493af0c008c0000263c000024",
INIT_15 => X"ac000000000000909090900003af27038f8f8fa30010a32414240010a3241000",
INIT_16 => X"a400009090a400009090ac00000000000090909090ac00000000000090909090",
INIT_17 => X"00008f9090a3a3af00000000000027909090909090a40300009090a400009090",
INIT_18 => X"afafafafafafafafaf002727032400100000009730143193241430932410a710",
INIT_19 => X"af2591242525258f919191242424242424242424242424242424242424afaf18",
INIT_1A => X"272726262693929292af000000000000242525252591919191ac000000000000",
INIT_1B => X"8f8f8f8f271400008faf000000000000262626262692929292ae000000000000",
INIT_1C => X"02021402020200028f2400142a020010020000afafafafaf2727038f8f8f8f8f",
INIT_1D => X"142497270c0214020c24000227afafafafafafafafafaf278f27038f8f8f8f8f",
INIT_1E => X"270202970200008f00029700240c028f2410001024100097241024142c009724",
INIT_1F => X"00008e8e0300100200008e8e000c028e27142c008e27272702af00100097020c",
INIT_20 => X"02140200008e8ea0140000249000028e8f001a0214248e0200278f2400142a00",
INIT_21 => X"8f8f8f8f8f8f8faf008f000c00000002029700020c02278f2614022626262797",
INIT_22 => X"278f00ac0324343c2703008f000caf3caf272703008f0000af278f27038f8f8f",
INIT_23 => X"0226ae30a002000c3c001a0000afafafafaf272703af8f008f8f020c0000afaf",
INIT_24 => X"0c243cac0c243424103cac0c24343c1030008c343caf2727038f8f8f8f8f0014",
INIT_25 => X"0024343c00ac2410002400ac343c343c00ac0c248fac0c24343c3c1400000c00",
INIT_26 => X"0000017f00ff202020202a0807070e0100000000000a00000000000000102410",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"00000084e00244e00200e042020000000062034202a560a4a01d8404a5059c1c",
INIT_01 => X"a086c6c5c406bb00bb00ba5a1abfb9b8afaeadacabaaa9a8a7a6a5a4a3a2a1bd",
INIT_02 => X"939291909b401bbd60bb60bbbabfb9b8afaeadacabaaa9a8a7a6a5a4a3a2a1a5",
INIT_03 => X"00e000c4e0000085a2e09f9d9c9e979695949392919002e09f9d9c9e97969594",
INIT_04 => X"a000b0b1b2bfbdbde000bf8400040000bfbd00e0004000828462420300400082",
INIT_05 => X"c543c686e30040420002e707080800a0bde0b0b1b2bf20504011100044508020",
INIT_06 => X"6263038440420042420242e042420240420062630302404200424202c0e00040",
INIT_07 => X"a062c505406303400042c2420240e04202424142026202630344e00200404200",
INIT_08 => X"6340424803c22e824800624a488a40e200a2c242020e2909c242028c0cc24202",
INIT_09 => X"0500a4a0a4a204a204bfbdbde000bf0500a4a0a4bfbd00e00040e5e720636361",
INIT_0A => X"4ac24343420203e002424142eb2c020a08080be7070c290960a00500bde000bf",
INIT_0B => X"e0c0a080b0b1b3b4b5bfb7b7b6b6b2b2bd62e002630300e00240c5c600438206",
INIT_0C => X"b0b1b2b3b4b5b6b7bf00006000a4e0e04000c0a0c04000802040000060005310",
INIT_0D => X"a6bfbdbde000bfa200a0a0a0bf84a2bdbde000bfa2000084a0a7a0bfa2bdbde0",
INIT_0E => X"00bfa000a00004a0bfbdbde000bfa000a00004a0bfbdbde000bf80004004a080",
INIT_0F => X"bde0454404430302b0bfa5a4a3a2a700a00004b0a700a00004b010b0bfbdbde0",
INIT_10 => X"000500a4060400050000041010b0bfbdbde04302bfa3a2a700a00004a202bfbd",
INIT_11 => X"10b0bfbdbde0b0bfa200000500a4060400050000041010b0bfbdbde0b0bfa200",
INIT_12 => X"024340000080620283400000bfbdbde0b0bfa200000500a40604000500000410",
INIT_13 => X"a0a0a082a20282020282020240438342824482b000b1bfbdbde000bf00008062",
INIT_14 => X"83428244820000a200a7425002a00004a0a0b11182a200a04250021010a00004",
INIT_15 => X"a24746064303028786838200e084bde0b0b1bf91000082028202000082024043",
INIT_16 => X"a362028382a362028382a247460643030287868382a247460643030287868382",
INIT_17 => X"8202858482a8a7a3666505620203bd888786858283a3e062028382a362028382",
INIT_18 => X"b0b1b2b3b4b5b6b7be00bdbde002020002430083824302830243e2830200a465",
INIT_19 => X"a80802e7294a6ba8234465898a8b8c8d8e8fd899909192d394959697dea4a5a0",
INIT_1A => X"18391031522203244502454404430302c68cadceef82a3c4e5c2454443020403",
INIT_1B => X"b5b6b7bede40e800a8c24544044303027394b5d6f782a3c4e562454404430302",
INIT_1C => X"2051403230004060821000400251804032c0a0b0b1b2b3bfbdbde0b0b1b2b3b4",
INIT_1D => X"6202a3a50000400000054000b0b0b1b2b3b4b5b6b7bebfbd82bde0b0b1b2b3bf",
INIT_1E => X"b10054a5804000820200a240050000a602000000026200a3020002404200a202",
INIT_1F => X"43002322c00060436440e4a3000040a6a4404200c2b6b5b720b0004000a22000",
INIT_20 => X"704042430023228340b082a563e56522a70000504707220040a4821000400252",
INIT_21 => X"b3b4b5b6b7bebf8300a3a60006c2024000a240400000b0a6d6408294b5f7dea2",
INIT_22 => X"bd848062e0026303bde000bf00008202bfbdbde000bf0040bfbd82bde0b0b1b2",
INIT_23 => X"1110424262700000128020a000b0b1b2b3bfbdbde082b050bf82000040a0b0bf",
INIT_24 => X"008404430003428400044300034202404200424202bfbdbde0b0b1b2b3bf0040",
INIT_25 => X"8363840400a06340c36300a7c606a5054062004283620002630305e040000000",
INIT_26 => X"0000024500ff00000000bc0406030c0200000000000d00000000000000006340",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"00000060006000002000001300000000040020000000ff180080130013009300",
INIT_01 => X"f8200000002000d800d800ff70000000000000000000000000000000000000ff",
INIT_02 => X"0000000060000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000201000000000000000000000000000000000000000000000000000",
INIT_04 => X"888000000000ff00000000130000000000ff000000ff00000000002000000000",
INIT_05 => X"100000100000000000000020002030000000000000001010ff10000000109000",
INIT_06 => X"000020000000000000200000000020ff000000002020000000000020100000ff",
INIT_07 => X"0000282838002040500010130000000020ffffff000000002000002000ff0000",
INIT_08 => X"ff40001000000000100000000010001000003013000000205813000020681300",
INIT_09 => X"00000030000012001400ff00000000000000300000ff000000ff10000000ffff",
INIT_0A => X"000000100010180000ffffff0000000000200000200000203000281800000000",
INIT_0B => X"a888a080000000000000000000000000ff0000000020000000ff100018001010",
INIT_0C => X"0000000000000000000001300100280030002820002801200028012020000000",
INIT_0D => X"0000ff000000000001000000000000ff00000000000138000000000000ff0000",
INIT_0E => X"000038013028000000ff0000000038013028000000ff00000000300128003810",
INIT_0F => X"0000101022101c16000000000000000130280000000130280000000000ff0000",
INIT_10 => X"010001000000010000000013000000ff000010120000000001302800000000ff",
INIT_11 => X"000000ff000000000000010001000000010000000013000000ff000000000000",
INIT_12 => X"00002000021000000020000200ff000000000000010001000000010000000013",
INIT_13 => X"0000008000008000000000000010000000008000020000ff0000000000021000",
INIT_14 => X"0000000080000200010000101030280000000000800001380010101300302800",
INIT_15 => X"00101032101c1600000000000080000000000080000080000000000080000010",
INIT_16 => X"0018120000001812000000101032101c160000000000101032101c1600000000",
INIT_17 => X"201280000000000018182a18141eff0000000000000000181200000018120000",
INIT_18 => X"00000000000000000038ff000000100010100080ff0000800000008000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"00000000000000000000101022101c160000000000000000000010101016221c",
INIT_1B => X"0000000000ff10000000101022101c1600000000000000000000101022101c16",
INIT_1C => X"1080ff108828f82080040000048098001090880000000000ff00000000000000",
INIT_1D => X"00000000022000200200f8200006060606060606060606f98000000000000000",
INIT_1E => X"0420900028f80080a12000900003200000000000000000000000000000000000",
INIT_1F => X"1000000088000018189000009803280000ff200000040404f006a00000003003",
INIT_20 => X"98ff101000000000ff102000001820000628009000000028f800800400000480",
INIT_21 => X"06060606060606801000300330303028200090280320000000ff100000000000",
INIT_22 => X"ff80100000000020000000000002800000ff0000000000f800ff800600060606",
INIT_23 => X"100000000018000020980088800000000000ff00008000100080300128800000",
INIT_24 => X"02110000040000110000000400002000000000002000ff0000000000000000ff",
INIT_25 => X"10008400180000ff1000180084000020380004ff800000000020200038000300",
INIT_26 => X"0000004c000100000000de020401000400000000000000000000000000ff00ff",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"00000000080044080000088000001100894c005c0004fd2a0000800080004301",
INIT_01 => X"0924504c400060125c1058fc0054504c4844403c3834302c2824201c18141098",
INIT_02 => X"0c080400000801681360115c5854504c4844403c3834302c2824201c18141000",
INIT_03 => X"00080c000810121900082c2824201c1814100c08040000082c2824201c181410",
INIT_04 => X"25251014181ce018080010288000008010e8000800fa00000100ff0000090000",
INIT_05 => X"2a00012100000808000004000800251120081014181c2521fb2a01d600212508",
INIT_06 => X"000800ff080100000800ff08000400fc080000080000080800000800250800f5",
INIT_07 => X"280007c025c8002525002144000008c000ffffff010002c00000080000fc0100",
INIT_08 => X"ff25ff04010000000700000100210324000021400001c000214c00c400214800",
INIT_09 => X"03f31025121103100318e02008001801f310251018e0000800e72a010001ffff",
INIT_0A => X"0407ff210142400000ffffff00000107c40001c0000fc8002521c02520080018",
INIT_0B => X"2525252510141c202430502c48285418c8000802c000000801eb2a01250021c3",
INIT_0C => X"1014181c2024282c30006a25444c250425f325250425352503252a2525e7ffff",
INIT_0D => X"1018e028080020106f1c181420ff38d828080020186f25ff1c14102038d83808",
INIT_0E => X"001825b02525041018e02008001825b02525061018e02008001825a225032525",
INIT_0F => X"280825210021000020241b1a19181aa22525651018a225258510022024d82008",
INIT_10 => X"6a01441007652a0400e7072c00181ce02808250020191818a22525b5100220d8",
INIT_11 => X"00181ce02008181c10006a0144100b652a0800e70b2c00181ce02008181c1000",
INIT_12 => X"80c0250026250ac0c025001010e82008181c10006a01441013652a1000e7132c",
INIT_13 => X"1814102720ff2702010280040525010140e02528522c30c81808001000102503",
INIT_14 => X"010140e02500521c6f2000218025256118141001271c6f250021802c00252506",
INIT_15 => X"002121002100001b1a19180008293808282c3027000227020480000827040425",
INIT_16 => X"0e21002d2c0c21002b2a0821210021000023222120042121002100001f1e1d1c",
INIT_17 => X"21002d1312050400212100210000f80504030201001208210031301021002f2e",
INIT_18 => X"080c1014181c20242825d008080380022b260033ff07ff32020cff3101100603",
INIT_19 => X"0020000120202000000000010203040506070408090a0b08101112130c00345b",
INIT_1A => X"1020202020000000000021210021000010202020200000000000212121000000",
INIT_1B => X"1c20242810ba2a00340021210021000010202020200000000000212100210000",
INIT_1C => X"2523f52a21250925290000020123250e2a25251014181c20d83008080c101418",
INIT_1D => X"79201c10b5257f25eb340925283034383c4044484c5054a82928081014181c20",
INIT_1E => X"2825211e2509002940251e2534872514086a006c070500200672280321001e05",
INIT_1F => X"21000c042500262b212500002587250028df000000302c3425282543001e2515",
INIT_20 => X"21dd2b21000c0400f72a21010021210828250b210d0100250928290000020123",
INIT_21 => X"3c4044484c50543525102187c0218025252225258725281810c42a011010101e",
INIT_22 => X"e839250008011000180800100068391810e818080010000910e8355808303438",
INIT_23 => X"2a0100ff002100c400250c25251014181c20d81808391021143925bd25251014",
INIT_24 => X"b27400004e5460b40700005866600008080000740010e828081014181c2000f7",
INIT_25 => X"2a017f1e250001fe2a0125007f1e6000250045ff110013ff6000000c2500a700",
INIT_26 => X"000008460000504c4440f0000000000002000100000000000000000000f101fe",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic
