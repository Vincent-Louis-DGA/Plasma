-------------------------------------------------------------------------------
-- Inferred BlockRAM with Initial Values
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Ram_Program is
  generic (
    N : integer := 4;                -- Width in bytes
    M : integer := 13);               -- Address width

  port (
    clk  : in  std_logic;
    wbe   : in  std_logic_vector(N-1 downto 0)   := (others => '0');
    addr : in  std_logic_vector(M-1 downto 0)   := (others => '0');
    din  : in  std_logic_vector(N*8-1 downto 0) := (others => '0');
    dout : out std_logic_vector(N*8-1 downto 0)
    );

end Ram_Program;

architecture logic of Ram_Program is

  type mem_file is array(0 to (2**M)-1) of std_logic_vector(N*8-1 downto 0);
  
  signal ram : mem_file := (
    -- Insert initial values below here, eg,
    -- 0 => X"0000",
    -- 1 => X"0001",
    -- <INIT_DATA>
0 => X"3C1C0001",1 => X"279C9F18",2 => X"3C050000",3 => X"24A51F58",
4 => X"3C040000",5 => X"24842060",6 => X"341D8000",7 => X"ACA00000",
8 => X"00A4182A",9 => X"1460FFFD",10 => X"24A50004",11 => X"3C020000",
12 => X"2442005C",13 => X"3C032000",14 => X"AC62004C",15 => X"0C0006DA",
16 => X"00000000",17 => X"08000011",18 => X"00000000",19 => X"3C020000",
20 => X"24422060",21 => X"03E00008",22 => X"00000000",23 => X"3C022000",
24 => X"03E00008",25 => X"AC440044",26 => X"40026000",27 => X"03E00008",
28 => X"40846000",29 => X"00000000",30 => X"00000000",31 => X"00000000",
32 => X"23BDFF98",33 => X"AFA10010",34 => X"AFA20014",35 => X"AFA30018",
36 => X"AFA4001C",37 => X"AFA50020",38 => X"AFA60024",39 => X"AFA70028",
40 => X"AFA8002C",41 => X"AFA90030",42 => X"AFAA0034",43 => X"AFAB0038",
44 => X"AFAC003C",45 => X"AFAD0040",46 => X"AFAE0044",47 => X"AFAF0048",
48 => X"AFB8004C",49 => X"AFB90050",50 => X"AFBF0054",51 => X"401A7000",
52 => X"235AFFFC",53 => X"AFBA0058",54 => X"0000D810",55 => X"AFBB005C",
56 => X"0000D812",57 => X"AFBB0060",58 => X"3C062000",59 => X"8CC40040",
60 => X"8CC5004C",61 => X"8CC60050",62 => X"00862024",63 => X"00A0F809",
64 => X"23A50000",65 => X"8FA10010",66 => X"8FA20014",67 => X"8FA30018",
68 => X"8FA4001C",69 => X"8FA50020",70 => X"8FA60024",71 => X"8FA70028",
72 => X"8FA8002C",73 => X"8FA90030",74 => X"8FAA0034",75 => X"8FAB0038",
76 => X"8FAC003C",77 => X"8FAD0040",78 => X"8FAE0044",79 => X"8FAF0048",
80 => X"8FB8004C",81 => X"8FB90050",82 => X"8FBF0054",83 => X"8FBA0058",
84 => X"8FBB005C",85 => X"03600011",86 => X"8FBB0060",87 => X"03600013",
88 => X"23BD0068",89 => X"341B0001",90 => X"03400008",91 => X"409B6000",
92 => X"AC900000",93 => X"AC910004",94 => X"AC920008",95 => X"AC93000C",
96 => X"AC940010",97 => X"AC950014",98 => X"AC960018",99 => X"AC97001C",
100 => X"AC9E0020",101 => X"AC9C0024",102 => X"AC9D0028",103 => X"AC9F002C",
104 => X"03E00008",105 => X"34020000",106 => X"8C900000",107 => X"8C910004",
108 => X"8C920008",109 => X"8C93000C",110 => X"8C940010",111 => X"8C950014",
112 => X"8C960018",113 => X"8C97001C",114 => X"8C9E0020",115 => X"8C9C0024",
116 => X"8C9D0028",117 => X"8C9F002C",118 => X"03E00008",119 => X"34A20000",
120 => X"00850019",121 => X"00001012",122 => X"00002010",123 => X"03E00008",
124 => X"ACC40000",125 => X"0000000C",126 => X"03E00008",127 => X"00000000",
128 => X"90820000",129 => X"00000000",130 => X"10400009",131 => X"00000000",
132 => X"3C032000",133 => X"304200FF",134 => X"AC620000",135 => X"24840001",
136 => X"90820000",137 => X"00000000",138 => X"1440FFFA",139 => X"00000000",
140 => X"03E00008",141 => X"00000000",142 => X"27BDFFE8",143 => X"AFBF0010",
144 => X"0C000080",145 => X"00000000",146 => X"3C040000",147 => X"0C000080",
148 => X"24841E44",149 => X"8FBF0010",150 => X"00000000",151 => X"03E00008",
152 => X"27BD0018",153 => X"27BDFFE0",154 => X"AFBF001C",155 => X"AFB20018",
156 => X"AFB10014",157 => X"AFB00010",158 => X"00008025",159 => X"00A08825",
160 => X"1A200008",161 => X"00809025",162 => X"02501021",163 => X"90440000",
164 => X"0C0000D6",165 => X"26100001",166 => X"0211102A",167 => X"1440FFFB",
168 => X"02501021",169 => X"02201025",170 => X"8FBF001C",171 => X"8FB20018",
172 => X"8FB10014",173 => X"8FB00010",174 => X"03E00008",175 => X"27BD0020",
176 => X"18A00011",177 => X"00003025",178 => X"3C082000",179 => X"35080008",
180 => X"3C072000",181 => X"34E70004",182 => X"8D020000",183 => X"00000000",
184 => X"30420008",185 => X"10400008",186 => X"00000000",187 => X"8CE30000",
188 => X"00861021",189 => X"24C60001",190 => X"A0430000",191 => X"00C5102A",
192 => X"1440FFF5",193 => X"00000000",194 => X"03E00008",195 => X"00C01025",
196 => X"3C022000",197 => X"34420008",198 => X"8C420000",199 => X"00000000",
200 => X"30420008",201 => X"14400008",202 => X"3C022000",203 => X"3C032000",
204 => X"34630008",205 => X"8C620000",206 => X"00000000",207 => X"30420008",
208 => X"1040FFFC",209 => X"3C022000",210 => X"34420004",211 => X"8C420000",
212 => X"03E00008",213 => X"304200FF",214 => X"3C022000",215 => X"34420008",
216 => X"8C420000",217 => X"00000000",218 => X"30420001",219 => X"10400008",
220 => X"308400FF",221 => X"3C032000",222 => X"34630008",223 => X"8C620000",
224 => X"00000000",225 => X"30420001",226 => X"1440FFFC",227 => X"00000000",
228 => X"3C022000",229 => X"03E00008",230 => X"AC440000",231 => X"18C0000E",
232 => X"00003825",233 => X"00871021",234 => X"90430000",235 => X"00A71021",
236 => X"90420000",237 => X"00000000",238 => X"14620007",239 => X"00000000",
240 => X"10600005",241 => X"00000000",242 => X"24E70001",243 => X"00E6102A",
244 => X"1440FFF5",245 => X"00871021",246 => X"10E60006",247 => X"00871021",
248 => X"90430000",249 => X"00A71021",250 => X"90420000",251 => X"10000002",
252 => X"00621023",253 => X"00001025",254 => X"03E00008",255 => X"00000000",
256 => X"90A20000",257 => X"00000000",258 => X"10400009",259 => X"00003025",
260 => X"90A20000",261 => X"24A50001",262 => X"00861821",263 => X"A0620000",
264 => X"90A20000",265 => X"00000000",266 => X"1440FFF9",267 => X"24C60001",
268 => X"00861021",269 => X"A0400000",270 => X"03E00008",271 => X"00C01025",
272 => X"00003825",273 => X"18A0000F",274 => X"00E03025",275 => X"00871021",
276 => X"90430000",277 => X"00000000",278 => X"2C62003A",279 => X"10400003",
280 => X"00061100",281 => X"10000002",282 => X"2442FFD0",283 => X"2442FFC9",
284 => X"00433021",285 => X"24E70001",286 => X"00E5102A",287 => X"1440FFF3",
288 => X"00000000",289 => X"03E00008",290 => X"00C01025",291 => X"00003025",
292 => X"18A0000A",293 => X"00C03825",294 => X"00861021",295 => X"90430000",
296 => X"24C60001",297 => X"00071040",298 => X"2442FFD0",299 => X"00433821",
300 => X"00C5102A",301 => X"1440FFF8",302 => X"00000000",303 => X"03E00008",
304 => X"00E01025",305 => X"00003825",306 => X"18A0000C",307 => X"00E03025",
308 => X"00871021",309 => X"90430000",310 => X"24E70001",311 => X"00061080",
312 => X"00461021",313 => X"00021040",314 => X"2442FFD0",315 => X"00433021",
316 => X"00E5102A",317 => X"1440FFF6",318 => X"00000000",319 => X"03E00008",
320 => X"00C01025",321 => X"27BDFFE8",322 => X"AFBF0010",323 => X"00A04825",
324 => X"AD200000",325 => X"90820000",326 => X"00002825",327 => X"10400012",
328 => X"24080064",329 => X"2442FFD0",330 => X"2C42000A",331 => X"14400009",
332 => X"00000000",333 => X"8D220000",334 => X"24840001",335 => X"24420001",
336 => X"AD220000",337 => X"90820000",338 => X"00000000",339 => X"1440FFF6",
340 => X"2442FFD0",341 => X"90820000",342 => X"00000000",343 => X"14400004",
344 => X"00851821",345 => X"AD200000",346 => X"1000003C",347 => X"00001025",
348 => X"90620000",349 => X"00000000",350 => X"10400022",351 => X"00000000",
352 => X"240C0001",353 => X"240B0078",354 => X"240A0062",355 => X"00603825",
356 => X"24A50001",357 => X"14AC000C",358 => X"24E70001",359 => X"90820001",
360 => X"00000000",361 => X"144B0003",362 => X"00000000",363 => X"10000010",
364 => X"24080078",365 => X"00000000",366 => X"144A0003",367 => X"00000000",
368 => X"1000000B",369 => X"24080062",370 => X"90E60000",371 => X"00000000",
372 => X"2CC30030",373 => X"24C2FFC6",374 => X"2C420007",375 => X"00621825",
376 => X"14600008",377 => X"2CC20047",378 => X"10400006",379 => X"00000000",
380 => X"90E20000",381 => X"00000000",382 => X"1440FFE6",383 => X"24A50001",
384 => X"24A5FFFF",385 => X"8D220000",386 => X"00000000",387 => X"00451021",
388 => X"AD220000",389 => X"24020078",390 => X"15020006",391 => X"24020062",
392 => X"24840002",393 => X"0C000110",394 => X"24A5FFFE",395 => X"1000000B",
396 => X"00000000",397 => X"00000000",398 => X"11020005",399 => X"00000000",
400 => X"0C000131",401 => X"00000000",402 => X"10000004",403 => X"00000000",
404 => X"24840002",405 => X"0C000123",406 => X"24A5FFFE",407 => X"8FBF0010",
408 => X"00000000",409 => X"03E00008",410 => X"27BD0018",411 => X"00A03825",
412 => X"24C2FFFE",413 => X"2C420023",414 => X"14400003",415 => X"00004025",
416 => X"1000002C",417 => X"A0A00000",418 => X"3C020000",419 => X"24491E48",
420 => X"00801825",421 => X"14C00002",422 => X"0086001A",423 => X"0007000D",
424 => X"2401FFFF",425 => X"14C10004",426 => X"3C018000",427 => X"14810002",
428 => X"00000000",429 => X"0006000D",430 => X"00002012",431 => X"00000000",
432 => X"00000000",433 => X"00860018",434 => X"00005812",435 => X"006B1023",
436 => X"00491021",437 => X"90420023",438 => X"25080001",439 => X"A0E20000",
440 => X"1480FFEB",441 => X"24E70001",442 => X"04610004",443 => X"2402002D",
444 => X"A0E20000",445 => X"24E70001",446 => X"25080001",447 => X"A0E00000",
448 => X"24E7FFFF",449 => X"00A7102B",450 => X"1040000A",451 => X"00000000",
452 => X"90A20000",453 => X"90E30000",454 => X"A0E20000",455 => X"A0A30000",
456 => X"24E7FFFF",457 => X"24A50001",458 => X"00A7102B",459 => X"1440FFF8",
460 => X"00000000",461 => X"03E00008",462 => X"01001025",463 => X"24020030",
464 => X"A0A20000",465 => X"24020078",466 => X"A0A20001",467 => X"24070002",
468 => X"2406001C",469 => X"2409000F",470 => X"3C020000",471 => X"24481E90",
472 => X"00C91804",473 => X"00831824",474 => X"00C31806",475 => X"306300FF",
476 => X"00681821",477 => X"90630000",478 => X"00A71021",479 => X"24E70001",
480 => X"24C6FFFC",481 => X"04C1FFF6",482 => X"A0430000",483 => X"00A71021",
484 => X"A0400000",485 => X"03E00008",486 => X"00E01025",487 => X"18C00016",
488 => X"00003825",489 => X"3C020000",490 => X"24491E90",491 => X"24A80001",
492 => X"00871821",493 => X"90620000",494 => X"00000000",495 => X"00021102",
496 => X"00491021",497 => X"90420000",498 => X"00000000",499 => X"A0A20000",
500 => X"90620000",501 => X"24E70001",502 => X"3042000F",503 => X"00491021",
504 => X"90420000",505 => X"24A50002",506 => X"A1020000",507 => X"00E6102A",
508 => X"1440FFEF",509 => X"25080002",510 => X"03E00008",511 => X"00000000",
512 => X"3C022000",513 => X"34420044",514 => X"AC440000",515 => X"8F828024",
516 => X"3C032000",517 => X"34630060",518 => X"24420001",519 => X"AF828024",
520 => X"03E00008",521 => X"AC620000",522 => X"27BDFFE8",523 => X"AFBF0010",
524 => X"3C022000",525 => X"34420060",526 => X"AC440000",527 => X"28822711",
528 => X"14400006",529 => X"00000000",530 => X"3C040000",531 => X"0C000080",
532 => X"24841EA4",533 => X"10000003",534 => X"00000000",535 => X"0C00020A",
536 => X"24840001",537 => X"8FBF0010",538 => X"00000000",539 => X"03E00008",
540 => X"27BD0018",541 => X"27BDFFE8",542 => X"AFBF0010",543 => X"0C000013",
544 => X"00000000",545 => X"AF828040",546 => X"00402825",547 => X"3C042000",
548 => X"34840060",549 => X"00051E03",550 => X"AC830000",551 => X"00051C03",
552 => X"AC830000",553 => X"00051A03",554 => X"AC830000",555 => X"AC850000",
556 => X"24050063",557 => X"2442018C",558 => X"AC450000",559 => X"24A5FFFF",
560 => X"04A1FFFD",561 => X"2442FFFC",562 => X"00002825",563 => X"3C032000",
564 => X"34630060",565 => X"AC650000",566 => X"24A50001",567 => X"28A20064",
568 => X"1440FFFC",569 => X"00000000",570 => X"8FBF0010",571 => X"00000000",
572 => X"03E00008",573 => X"27BD0018",574 => X"27BDFFD8",575 => X"AFBF0024",
576 => X"AFB20020",577 => X"AFB1001C",578 => X"AFB00018",579 => X"00808825",
580 => X"0C000141",581 => X"27A50010",582 => X"8FB00010",583 => X"00409025",
584 => X"27A50010",585 => X"0C000141",586 => X"02302021",587 => X"00121A00",
588 => X"00629021",589 => X"8FA20010",590 => X"27A50010",591 => X"02028021",
592 => X"0C000141",593 => X"02302021",594 => X"00121A00",595 => X"00629021",
596 => X"8FA20010",597 => X"27A50010",598 => X"02028021",599 => X"0C000141",
600 => X"02302021",601 => X"8FBF0024",602 => X"00121A00",603 => X"8FB20020",
604 => X"8FB1001C",605 => X"8FB00018",606 => X"00621021",607 => X"03E00008",
608 => X"27BD0028",609 => X"27BDFFE0",610 => X"AFBF0018",611 => X"AFB10014",
612 => X"AFB00010",613 => X"AFA40020",614 => X"27A40020",615 => X"00A08025",
616 => X"0C0001E7",617 => X"24060001",618 => X"2411002E",619 => X"A2110002",
620 => X"27A40021",621 => X"26050003",622 => X"0C0001E7",623 => X"24060001",
624 => X"A2110005",625 => X"27A40022",626 => X"26050006",627 => X"0C0001E7",
628 => X"24060001",629 => X"A2110008",630 => X"27A40023",631 => X"26050009",
632 => X"0C0001E7",633 => X"24060001",634 => X"8FBF0018",635 => X"8FB10014",
636 => X"8FB00010",637 => X"03E00008",638 => X"27BD0020",639 => X"27BDFFC8",
640 => X"AFBF0034",641 => X"AFBE0030",642 => X"AFB7002C",643 => X"AFB60028",
644 => X"AFB50024",645 => X"AFB40020",646 => X"AFB3001C",647 => X"AFB20018",
648 => X"AFB10014",649 => X"AFB00010",650 => X"AFA40038",651 => X"00008025",
652 => X"3C112001",653 => X"36315020",654 => X"3C142001",655 => X"36944000",
656 => X"3C132001",657 => X"36735030",658 => X"241E0800",659 => X"24170806",
660 => X"3C16F000",661 => X"3C154000",662 => X"3C120001",663 => X"36520800",
664 => X"02111026",665 => X"8C420000",666 => X"00000000",667 => X"3042FFFF",
668 => X"10400017",669 => X"02131026",670 => X"8C420000",671 => X"02142026",
672 => X"3042FFFF",673 => X"105E000A",674 => X"00401825",675 => X"1057000E",
676 => X"2C620600",677 => X"1040000F",678 => X"02111026",679 => X"8C830000",
680 => X"00000000",681 => X"00761024",682 => X"14550005",683 => X"00000000",
684 => X"0C000722",685 => X"00000000",686 => X"10000006",687 => X"02111026",
688 => X"14720004",689 => X"02111026",690 => X"0C00045D",691 => X"02002825",
692 => X"02111026",693 => X"AC400000",694 => X"26100800",695 => X"2E020801",
696 => X"1440FFE0",697 => X"02111026",698 => X"8F828018",699 => X"8FA60038",
700 => X"00000000",701 => X"AC460000",702 => X"8FBF0034",703 => X"8FBE0030",
704 => X"8FB7002C",705 => X"8FB60028",706 => X"8FB50024",707 => X"8FB40020",
708 => X"8FB3001C",709 => X"8FB20018",710 => X"8FB10014",711 => X"8FB00010",
712 => X"03E00008",713 => X"27BD0038",714 => X"3C022001",715 => X"34420024",
716 => X"3084FFFF",717 => X"AC440000",718 => X"3C022001",719 => X"34420028",
720 => X"30A5FFFF",721 => X"AC450000",722 => X"3C022001",723 => X"3442002C",
724 => X"30C6FFFF",725 => X"AC460000",726 => X"3C022001",727 => X"34425020",
728 => X"AC400000",729 => X"3C022001",730 => X"34425820",731 => X"03E00008",
732 => X"AC400000",733 => X"8F83801C",734 => X"27BDFFE8",735 => X"AFBF0010",
736 => X"3C020000",737 => X"244209FC",738 => X"AC620000",739 => X"8F838020",
740 => X"24020004",741 => X"AC620000",742 => X"8F828014",743 => X"24040001",
744 => X"0C00001A",745 => X"AC400000",746 => X"8FBF0010",747 => X"00000000",
748 => X"03E00008",749 => X"27BD0018",750 => X"00001825",751 => X"30A5FFFF",
752 => X"10A00008",753 => X"00603025",754 => X"94820000",755 => X"24630002",
756 => X"3063FFFF",757 => X"00C23021",758 => X"0065102B",759 => X"1440FFFA",
760 => X"24840002",761 => X"30C3FFFF",762 => X"00061402",763 => X"00623021",
764 => X"00061027",765 => X"03E00008",766 => X"3042FFFF",767 => X"3C022001",
768 => X"34423024",769 => X"3084FFFF",770 => X"AC440000",771 => X"3C022001",
772 => X"34423028",773 => X"30A5FFFF",774 => X"AC450000",775 => X"3C022001",
776 => X"3442302C",777 => X"30C6FFFF",778 => X"03E00008",779 => X"AC460000",
780 => X"3C022001",781 => X"34423000",782 => X"8C420000",783 => X"00000000",
784 => X"30420004",785 => X"10400008",786 => X"00000000",787 => X"3C032001",
788 => X"34633000",789 => X"8C620000",790 => X"00000000",791 => X"30420004",
792 => X"1440FFFC",793 => X"00000000",794 => X"03E00008",795 => X"00000000",
796 => X"3C022001",797 => X"34423000",798 => X"8C420000",799 => X"00000000",
800 => X"30420004",801 => X"10400007",802 => X"3C032001",803 => X"34633000",
804 => X"8C620000",805 => X"00000000",806 => X"30420004",807 => X"1440FFFC",
808 => X"00000000",809 => X"3C022001",810 => X"34423020",811 => X"AC440000",
812 => X"3C032001",813 => X"34633000",814 => X"24020002",815 => X"03E00008",
816 => X"AC620000",817 => X"8C820010",818 => X"00000000",819 => X"ACA20004",
820 => X"8C82000C",821 => X"00000000",822 => X"ACA20000",823 => X"90820009",
824 => X"03E00008",825 => X"A0A20008",826 => X"8C820004",827 => X"00000000",
828 => X"ACA20004",829 => X"8C820000",830 => X"00000000",831 => X"ACA20000",
832 => X"90820008",833 => X"03E00008",834 => X"A0A20008",835 => X"8CA30000",
836 => X"00000000",837 => X"10600005",838 => X"00000000",839 => X"8C820000",
840 => X"00000000",841 => X"14620012",842 => X"00001025",843 => X"8CA30004",
844 => X"00000000",845 => X"10600005",846 => X"00000000",847 => X"8C820004",
848 => X"00000000",849 => X"1462000A",850 => X"00001025",851 => X"90A50008",
852 => X"00000000",853 => X"10A00006",854 => X"24020001",855 => X"90830008",
856 => X"00000000",857 => X"14A30002",858 => X"00001025",859 => X"24020001",
860 => X"03E00008",861 => X"00000000",862 => X"27BDFFC8",863 => X"AFBF0030",
864 => X"AFB5002C",865 => X"AFB40028",866 => X"AFB30024",867 => X"AFB20020",
868 => X"AFB1001C",869 => X"AFB00018",870 => X"00808825",871 => X"3C040000",
872 => X"24841EB0",873 => X"0C000099",874 => X"24050002",875 => X"3C020000",
876 => X"24501F60",877 => X"8E220020",878 => X"27A40010",879 => X"02002825",
880 => X"24060004",881 => X"0C0001E7",882 => X"AFA20010",883 => X"02002025",
884 => X"0C000099",885 => X"24050008",886 => X"0C0000D6",887 => X"2404003B",
888 => X"8FA30010",889 => X"8F828044",890 => X"00000000",891 => X"14620053",
892 => X"02002825",893 => X"8E24002C",894 => X"0C000261",895 => X"AFA40010",
896 => X"02002025",897 => X"0C000099",898 => X"2405000B",899 => X"0C0000D6",
900 => X"2404003B",901 => X"93828030",902 => X"00000000",903 => X"14400004",
904 => X"00000000",905 => X"8FA20010",906 => X"00000000",907 => X"AF82802C",
908 => X"8E240030",909 => X"02002825",910 => X"0C000261",911 => X"AFA40010",
912 => X"02002025",913 => X"0C000099",914 => X"2405000B",915 => X"0C0000D6",
916 => X"2404003B",917 => X"93828030",918 => X"00000000",919 => X"14400004",
920 => X"00000000",921 => X"8FA20010",922 => X"00000000",923 => X"AF828034",
924 => X"2631010C",925 => X"00009025",926 => X"241500FF",927 => X"24140001",
928 => X"02009825",929 => X"92230000",930 => X"00000000",931 => X"1075002B",
932 => X"00000000",933 => X"92300001",934 => X"00000000",935 => X"2E020020",
936 => X"10400026",937 => X"38630033",938 => X"2C630001",939 => X"3A020004",
940 => X"2C420001",941 => X"00621824",942 => X"10600010",943 => X"00000000",
944 => X"93828030",945 => X"00000000",946 => X"1454000C",947 => X"00000000",
948 => X"92220002",949 => X"92230003",950 => X"92240004",951 => X"92250005",
952 => X"00021600",953 => X"00031C00",954 => X"00431021",955 => X"00042200",
956 => X"00441021",957 => X"00451021",958 => X"AF828028",959 => X"02202025",
960 => X"02602825",961 => X"0C0001E7",962 => X"26060002",963 => X"02602025",
964 => X"00102840",965 => X"0C000099",966 => X"24A50004",967 => X"0C0000D6",
968 => X"2404003B",969 => X"02301021",970 => X"24510002",971 => X"26520001",
972 => X"2A42000A",973 => X"1440FFD3",974 => X"00000000",975 => X"8FBF0030",
976 => X"8FB5002C",977 => X"8FB40028",978 => X"8FB30024",979 => X"8FB20020",
980 => X"8FB1001C",981 => X"8FB00018",982 => X"03E00008",983 => X"27BD0038",
984 => X"27BDFFE0",985 => X"AFBF0018",986 => X"AFB10014",987 => X"AFB00010",
988 => X"00808025",989 => X"3C040000",990 => X"24841EB4",991 => X"00A08825",
992 => X"0C000099",993 => X"24050002",994 => X"26040014",995 => X"3C100000",
996 => X"26101F60",997 => X"02002825",998 => X"0C0001E7",999 => X"24060002",
1000 => X"02002025",1001 => X"0C000099",1002 => X"24050004",1003 => X"0C0000D6",
1004 => X"2404003B",1005 => X"8F838038",1006 => X"24020003",1007 => X"10620010",
1008 => X"00000000",1009 => X"8F828038",1010 => X"02202025",1011 => X"3C100000",
1012 => X"24420001",1013 => X"AF828038",1014 => X"8F858038",1015 => X"26101FE0",
1016 => X"00052940",1017 => X"0C00033A",1018 => X"00B02821",1019 => X"8F828038",
1020 => X"00000000",1021 => X"00021140",1022 => X"00501021",1023 => X"AC40001C",
1024 => X"8FBF0018",1025 => X"8FB10014",1026 => X"8FB00010",1027 => X"03E00008",
1028 => X"27BD0020",1029 => X"27BDFFE8",1030 => X"AFBF0014",1031 => X"AFB00010",
1032 => X"00808025",1033 => X"0C0000D6",1034 => X"24040054",1035 => X"26040014",
1036 => X"3C100000",1037 => X"26101F60",1038 => X"02002825",1039 => X"0C0001E7",
1040 => X"24060002",1041 => X"02002025",1042 => X"0C000099",1043 => X"24050004",
1044 => X"0C0000D6",1045 => X"2404003B",1046 => X"8FBF0014",1047 => X"8FB00010",
1048 => X"03E00008",1049 => X"27BD0018",1050 => X"27BDFFD8",1051 => X"AFBF0020",
1052 => X"AFB1001C",1053 => X"AFB00018",1054 => X"00808825",1055 => X"96220014",
1056 => X"96230016",1057 => X"3C040000",1058 => X"24841EB8",1059 => X"24050002",
1060 => X"A7A20010",1061 => X"0C000099",1062 => X"A7A30012",1063 => X"27A40010",
1064 => X"3C100000",1065 => X"26101F60",1066 => X"02002825",1067 => X"0C0001E7",
1068 => X"24060002",1069 => X"02002025",1070 => X"0C000099",1071 => X"24050004",
1072 => X"0C0000D6",1073 => X"2404003B",1074 => X"27A40012",1075 => X"02002825",
1076 => X"0C0001E7",1077 => X"24060002",1078 => X"02002025",1079 => X"0C000099",
1080 => X"24050004",1081 => X"0C0000D6",1082 => X"2404003B",1083 => X"97A30012",
1084 => X"24020044",1085 => X"14620003",1086 => X"00000000",1087 => X"0C00035E",
1088 => X"02202025",1089 => X"8FBF0020",1090 => X"8FB1001C",1091 => X"8FB00018",
1092 => X"03E00008",1093 => X"27BD0028",1094 => X"27BDFFE8",1095 => X"AFBF0014",
1096 => X"AFB00010",1097 => X"00808025",1098 => X"3C040000",1099 => X"24841EBC",
1100 => X"0C000099",1101 => X"24050002",1102 => X"26040014",1103 => X"3C100000",
1104 => X"26101F60",1105 => X"02002825",1106 => X"0C0001E7",1107 => X"24060002",
1108 => X"02002025",1109 => X"0C000099",1110 => X"24050004",1111 => X"0C0000D6",
1112 => X"2404003B",1113 => X"8FBF0014",1114 => X"8FB00010",1115 => X"03E00008",
1116 => X"27BD0018",1117 => X"27BDFFE8",1118 => X"AFBF0014",1119 => X"AFB00010",
1120 => X"00A08025",1121 => X"3C040000",1122 => X"24841EC0",1123 => X"0C000099",
1124 => X"24050002",1125 => X"8F838038",1126 => X"24020003",1127 => X"10620023",
1128 => X"00000000",1129 => X"8F828038",1130 => X"3C052001",1131 => X"34A55034",
1132 => X"3C062001",1133 => X"34C65038",1134 => X"3C072001",1135 => X"34E7503C",
1136 => X"3C040000",1137 => X"24841FE0",1138 => X"24030001",1139 => X"02052826",
1140 => X"02063026",1141 => X"24420001",1142 => X"AF828038",1143 => X"8F828038",
1144 => X"02073826",1145 => X"00021140",1146 => X"00441021",1147 => X"AC43001C",
1148 => X"8F828038",1149 => X"8CA30000",1150 => X"00021140",1151 => X"00441021",
1152 => X"AC43000C",1153 => X"8F828038",1154 => X"8CC30000",1155 => X"00021140",
1156 => X"00441021",1157 => X"AC430010",1158 => X"8F828038",1159 => X"8CE30000",
1160 => X"00021140",1161 => X"00441021",1162 => X"AC430014",1163 => X"8FBF0014",
1164 => X"8FB00010",1165 => X"03E00008",1166 => X"27BD0018",1167 => X"27BDFFE8",
1168 => X"AFBF0014",1169 => X"AFB00010",1170 => X"24024500",1171 => X"3C012001",
1172 => X"A4222000",1173 => X"3C012001",1174 => X"A4242002",1175 => X"3C026DF3",
1176 => X"3C012001",1177 => X"AC222004",1178 => X"30A580FF",1179 => X"34A58000",
1180 => X"3C012001",1181 => X"A4252008",1182 => X"3C102001",1183 => X"3610200A",
1184 => X"A6000000",1185 => X"3C012001",1186 => X"AC26200C",1187 => X"3C012001",
1188 => X"AC272010",1189 => X"3C042001",1190 => X"34842000",1191 => X"0C0002EE",
1192 => X"24050014",1193 => X"A6020000",1194 => X"8FBF0014",1195 => X"8FB00010",
1196 => X"03E00008",1197 => X"27BD0018",1198 => X"27BDFFE0",1199 => X"AFBF0018",
1200 => X"AFB10014",1201 => X"AFB00010",1202 => X"00801825",1203 => X"00C08825",
1204 => X"3224FFFF",1205 => X"00A01025",1206 => X"24050001",1207 => X"00E08025",
1208 => X"3210FFFF",1209 => X"00603025",1210 => X"0C00048F",1211 => X"00403825",
1212 => X"24020800",1213 => X"3C012001",1214 => X"A4222014",1215 => X"3C012001",
1216 => X"A4202016",1217 => X"24020001",1218 => X"3C012001",1219 => X"A4222018",
1220 => X"3C012001",1221 => X"A430201A",1222 => X"3C042001",1223 => X"3484201C",
1224 => X"2625FFE4",1225 => X"18A00008",1226 => X"00001825",1227 => X"3062000F",
1228 => X"24420061",1229 => X"A0820000",1230 => X"24630001",1231 => X"0065102A",
1232 => X"1440FFFA",1233 => X"24840001",1234 => X"3C042001",1235 => X"34842014",
1236 => X"2625FFEC",1237 => X"0C0002EE",1238 => X"30A5FFFF",1239 => X"8FBF0018",
1240 => X"8FB10014",1241 => X"8FB00010",1242 => X"3C012001",1243 => X"A4222016",
1244 => X"03E00008",1245 => X"27BD0020",1246 => X"27BDFFD8",1247 => X"AFB20018",
1248 => X"8FB20038",1249 => X"AFBF0024",1250 => X"AFB40020",1251 => X"AFB3001C",
1252 => X"AFB10014",1253 => X"AFB00010",1254 => X"3C132001",1255 => X"36732014",
1256 => X"00801025",1257 => X"00A01825",1258 => X"00C08025",1259 => X"00E08825",
1260 => X"3210FFFF",1261 => X"3231FFFF",1262 => X"24050011",1263 => X"00403025",
1264 => X"00603825",1265 => X"2654001C",1266 => X"0C00048F",1267 => X"3284FFFF",
1268 => X"A6700000",1269 => X"A6710002",1270 => X"26520008",1271 => X"A6720004",
1272 => X"A6600006",1273 => X"8FBF0024",1274 => X"02801025",1275 => X"8FB40020",
1276 => X"8FB3001C",1277 => X"8FB20018",1278 => X"8FB10014",1279 => X"8FB00010",
1280 => X"03E00008",1281 => X"27BD0028",1282 => X"27BDFFE0",1283 => X"AFBF001C",
1284 => X"AFB00018",1285 => X"00808025",1286 => X"3404FFFF",1287 => X"00802825",
1288 => X"0C0002FF",1289 => X"00803025",1290 => X"3C052001",1291 => X"34A5201C",
1292 => X"3C020101",1293 => X"34420600",1294 => X"ACA20000",1295 => X"3C012001",
1296 => X"AC302020",1297 => X"3C012001",1298 => X"AC202024",1299 => X"3C012001",
1300 => X"AC202028",1301 => X"3C012001",1302 => X"AC20202C",1303 => X"3C012001",
1304 => X"AC202030",1305 => X"3C012001",1306 => X"AC202034",1307 => X"2402020A",
1308 => X"3C012001",1309 => X"A4222038",1310 => X"24023544",1311 => X"3C012001",
1312 => X"A422203A",1313 => X"24025441",1314 => X"3C012001",1315 => X"A422203C",
1316 => X"24030022",1317 => X"240400C9",1318 => X"00A31021",1319 => X"A0400000",
1320 => X"2484FFFF",1321 => X"0481FFFC",1322 => X"24630001",1323 => X"3C026382",
1324 => X"34425363",1325 => X"ACA200EC",1326 => X"24023501",1327 => X"A4A200F0",
1328 => X"24020001",1329 => X"A0A200F2",1330 => X"240200FF",1331 => X"A0A200F3",
1332 => X"240300F4",1333 => X"AFA30010",1334 => X"00002025",1335 => X"2405FFFF",
1336 => X"24060044",1337 => X"0C0004DE",1338 => X"24070043",1339 => X"8FBF001C",
1340 => X"8FB00018",1341 => X"03E00008",1342 => X"27BD0020",1343 => X"8F838034",
1344 => X"3C023501",1345 => X"34420300",1346 => X"3C012001",1347 => X"AC22210C",
1348 => X"24023204",1349 => X"3C012001",1350 => X"A4222110",1351 => X"240200FF",
1352 => X"3C012001",1353 => X"A0222116",1354 => X"27BDFFE0",1355 => X"240200FB",
1356 => X"AFA20010",1357 => X"8F82802C",1358 => X"AFBF0018",1359 => X"00002025",
1360 => X"2405FFFF",1361 => X"24060044",1362 => X"24070043",1363 => X"3C012001",
1364 => X"AC232030",1365 => X"8F83802C",1366 => X"00021402",1367 => X"3C012001",
1368 => X"A4222112",1369 => X"3C012001",1370 => X"0C0004DE",1371 => X"A4232114",
1372 => X"8FBF0018",1373 => X"00000000",1374 => X"03E00008",1375 => X"27BD0020",
1376 => X"27BDFFD8",1377 => X"AFBF0024",1378 => X"AFB40020",1379 => X"AFB3001C",
1380 => X"AFB20018",1381 => X"AFB10014",1382 => X"AFB00010",1383 => X"3C020000",
1384 => X"24431F1C",1385 => X"AC600004",1386 => X"AC401F1C",1387 => X"24020011",
1388 => X"A0620008",1389 => X"3C023544",1390 => X"34425441",1391 => X"AF828044",
1392 => X"00009825",1393 => X"3C102001",1394 => X"36103000",1395 => X"3C142001",
1396 => X"36943020",1397 => X"24120002",1398 => X"8F82802C",1399 => X"00000000",
1400 => X"14400038",1401 => X"00008825",1402 => X"AF80802C",1403 => X"A3808030",
1404 => X"AF808028",1405 => X"8E020000",1406 => X"00000000",1407 => X"30420004",
1408 => X"10400007",1409 => X"3C032001",1410 => X"34633000",1411 => X"8C620000",
1412 => X"00000000",1413 => X"30420004",1414 => X"1440FFFC",1415 => X"00000000",
1416 => X"8F828044",1417 => X"00000000",1418 => X"24420001",1419 => X"AF828044",
1420 => X"8F848044",1421 => X"0C000502",1422 => X"00000000",1423 => X"AE820000",
1424 => X"AE120000",1425 => X"8E020000",1426 => X"00000000",1427 => X"30420004",
1428 => X"10400007",1429 => X"3C032001",1430 => X"34633000",1431 => X"8C620000",
1432 => X"00000000",1433 => X"30420004",1434 => X"1440FFFC",1435 => X"00000000",
1436 => X"00001825",1437 => X"2402270F",1438 => X"2442FFFF",1439 => X"0441FFFF",
1440 => X"2442FFFF",1441 => X"8F82802C",1442 => X"00000000",1443 => X"14400005",
1444 => X"00000000",1445 => X"24630001",1446 => X"286203E8",1447 => X"1440FFF6",
1448 => X"2402270F",1449 => X"26310001",1450 => X"2A22000A",1451 => X"10400006",
1452 => X"24020001",1453 => X"8F82802C",1454 => X"00000000",1455 => X"1040FFCA",
1456 => X"00000000",1457 => X"24020001",1458 => X"A3828030",1459 => X"8E020000",
1460 => X"00000000",1461 => X"30420004",1462 => X"10400007",1463 => X"3C032001",
1464 => X"34633000",1465 => X"8C620000",1466 => X"00000000",1467 => X"30420004",
1468 => X"1440FFFC",1469 => X"00000000",1470 => X"0C00053F",1471 => X"00000000",
1472 => X"AE820000",1473 => X"AE120000",1474 => X"8E020000",1475 => X"00000000",
1476 => X"30420004",1477 => X"10400007",1478 => X"3C032001",1479 => X"34633000",
1480 => X"8C620000",1481 => X"00000000",1482 => X"30420004",1483 => X"1440FFFC",
1484 => X"00000000",1485 => X"00001825",1486 => X"2402270F",1487 => X"2442FFFF",
1488 => X"0441FFFF",1489 => X"2442FFFF",1490 => X"8F828028",1491 => X"00000000",
1492 => X"10400004",1493 => X"00000000",1494 => X"A3928030",1495 => X"10000009",
1496 => X"00000000",1497 => X"24630001",1498 => X"286203E8",1499 => X"1440FFF3",
1500 => X"2402270F",1501 => X"26730001",1502 => X"2A62000A",1503 => X"1440FF96",
1504 => X"00000000",1505 => X"8FBF0024",1506 => X"8FB40020",1507 => X"8FB3001C",
1508 => X"8FB20018",1509 => X"8FB10014",1510 => X"8FB00010",1511 => X"03E00008",
1512 => X"27BD0028",1513 => X"8F82802C",1514 => X"27BDFFD8",1515 => X"AFBF0020",
1516 => X"AFB3001C",1517 => X"AFB20018",1518 => X"AFB10014",1519 => X"AFB00010",
1520 => X"00E09825",1521 => X"3090FFFF",1522 => X"30B1FFFF",1523 => X"1040003C",
1524 => X"30D2FFFF",1525 => X"0C00030C",1526 => X"00000000",1527 => X"02002025",
1528 => X"02202825",1529 => X"0C0002FF",1530 => X"02403025",1531 => X"3C102001",
1532 => X"36103030",1533 => X"24020806",1534 => X"AE020000",1535 => X"24020001",
1536 => X"3C012001",1537 => X"A4222000",1538 => X"24020800",1539 => X"3C012001",
1540 => X"A4222002",1541 => X"24020604",1542 => X"3C012001",1543 => X"A4222004",
1544 => X"24020002",1545 => X"3C012001",1546 => X"A4222006",1547 => X"3C012001",
1548 => X"A4202012",1549 => X"3C012001",1550 => X"A4202014",1551 => X"3C012001",
1552 => X"A4202016",1553 => X"00131402",1554 => X"3C012001",1555 => X"A4222018",
1556 => X"3C012001",1557 => X"A433201A",1558 => X"3C032001",1559 => X"34630024",
1560 => X"8C630000",1561 => X"3C042001",1562 => X"34840028",1563 => X"8C850000",
1564 => X"3C022001",1565 => X"3442002C",1566 => X"8C420000",1567 => X"3C012001",
1568 => X"A422200C",1569 => X"8F82802C",1570 => X"3C012001",1571 => X"A4232008",
1572 => X"8F83802C",1573 => X"3C012001",1574 => X"A425200A",1575 => X"00021402",
1576 => X"3C012001",1577 => X"A422200E",1578 => X"3C012001",1579 => X"A4232010",
1580 => X"0C00031C",1581 => X"2404002E",1582 => X"24020800",1583 => X"AE020000",
1584 => X"8FBF0020",1585 => X"8FB3001C",1586 => X"8FB20018",1587 => X"8FB10014",
1588 => X"8FB00010",1589 => X"03E00008",1590 => X"27BD0028",1591 => X"27BDFFD8",
1592 => X"AFB3001C",1593 => X"8F938038",1594 => X"24020004",1595 => X"AFBF0020",
1596 => X"AFB20018",1597 => X"AFB10014",1598 => X"AFB00010",1599 => X"AF828038",
1600 => X"06600036",1601 => X"2402FFFF",1602 => X"3C020000",1603 => X"24421FE0",
1604 => X"00131940",1605 => X"00622021",1606 => X"8C83001C",1607 => X"24020001",
1608 => X"14620004",1609 => X"00000000",1610 => X"3C040000",1611 => X"10000007",
1612 => X"24841EC8",1613 => X"8C82001C",1614 => X"00000000",1615 => X"14400005",
1616 => X"00000000",1617 => X"3C040000",1618 => X"24841ECC",1619 => X"0C000099",
1620 => X"24050001",1621 => X"26640030",1622 => X"0C0000D6",1623 => X"308400FF",
1624 => X"0C0000D6",1625 => X"2404000A",1626 => X"3C042001",1627 => X"34843024",
1628 => X"8C900000",1629 => X"3C032001",1630 => X"34633028",1631 => X"8C710000",
1632 => X"3C022001",1633 => X"3442302C",1634 => X"8C520000",1635 => X"3C020000",
1636 => X"24421FE0",1637 => X"00131940",1638 => X"00621821",1639 => X"8C64000C",
1640 => X"8C650010",1641 => X"8C660014",1642 => X"8C670018",1643 => X"3084FFFF",
1644 => X"30A5FFFF",1645 => X"30C6FFFF",1646 => X"3210FFFF",1647 => X"3231FFFF",
1648 => X"0C0005E9",1649 => X"3252FFFF",1650 => X"02002025",1651 => X"02202825",
1652 => X"0C0002FF",1653 => X"02403025",1654 => X"2662FFFF",1655 => X"AF828038",
1656 => X"8FBF0020",1657 => X"8FB3001C",1658 => X"8FB20018",1659 => X"8FB10014",
1660 => X"8FB00010",1661 => X"03E00008",1662 => X"27BD0028",1663 => X"27BDFFD0",
1664 => X"AFBF002C",1665 => X"AFB40028",1666 => X"AFB30024",1667 => X"AFB20020",
1668 => X"AFB1001C",1669 => X"AFB00018",1670 => X"2404020A",1671 => X"24053544",
1672 => X"0C0002CA",1673 => X"24065441",1674 => X"0C000560",1675 => X"00000000",
1676 => X"3C040000",1677 => X"24841ED0",1678 => X"0C000099",1679 => X"2405000D",
1680 => X"8F84802C",1681 => X"3C100000",1682 => X"26101FA0",1683 => X"02002825",
1684 => X"00009025",1685 => X"0C000261",1686 => X"3414EA60",1687 => X"02002025",
1688 => X"0C000099",1689 => X"2405000B",1690 => X"3C040000",1691 => X"24841EE0",
1692 => X"0C000099",1693 => X"24050001",1694 => X"3C040000",1695 => X"24841EE4",
1696 => X"0C000099",1697 => X"24050007",1698 => X"27848028",1699 => X"02002825",
1700 => X"0C0001E7",1701 => X"24060004",1702 => X"02002025",1703 => X"0C000099",
1704 => X"24050008",1705 => X"0C0000D6",1706 => X"2404000A",1707 => X"8F87802C",
1708 => X"3404FFFF",1709 => X"00802825",1710 => X"0C0005E9",1711 => X"00803025",
1712 => X"240470F3",1713 => X"34059500",1714 => X"0C0002FF",1715 => X"2406721F",
1716 => X"3C040000",1717 => X"0C00023E",1718 => X"24841EEC",1719 => X"3C030000",
1720 => X"24641F1C",1721 => X"A0800008",1722 => X"AC601F1C",1723 => X"8F83802C",
1724 => X"00409825",1725 => X"AC830004",1726 => X"0C000637",1727 => X"24110400",
1728 => X"0C00030C",1729 => X"3C102001",1730 => X"3610201C",1731 => X"00001825",
1732 => X"A2030000",1733 => X"24630001",1734 => X"0071102A",1735 => X"1440FFFC",
1736 => X"26100001",1737 => X"8F84802C",1738 => X"AFB10010",1739 => X"02602825",
1740 => X"00003025",1741 => X"02543821",1742 => X"30E7FFFF",1743 => X"0C0004DE",
1744 => X"26520001",1745 => X"0C00031C",1746 => X"00402025",1747 => X"2E420020",
1748 => X"1440FFE9",1749 => X"00000000",1750 => X"0C000637",1751 => X"00000000",
1752 => X"1000FFFD",1753 => X"00000000",1754 => X"27BDFFA0",1755 => X"AFBF0058",
1756 => X"AFB10054",1757 => X"AFB00050",1758 => X"3C020123",1759 => X"34424567",
1760 => X"AC020010",1761 => X"3C040000",1762 => X"0C000080",1763 => X"24841EFC",
1764 => X"0C00067F",1765 => X"00000000",1766 => X"0C00021D",1767 => X"00000000",
1768 => X"0C00020A",1769 => X"00002025",1770 => X"00000000",1771 => X"00000000",
1772 => X"00000000",1773 => X"00000000",1774 => X"00000000",1775 => X"00000000",
1776 => X"00000000",1777 => X"00000000",1778 => X"3C022000",1779 => X"34420070",
1780 => X"8C510000",1781 => X"3C102000",1782 => X"36100060",1783 => X"26310001",
1784 => X"AE110000",1785 => X"00000000",1786 => X"00000000",1787 => X"00000000",
1788 => X"00000000",1789 => X"00000000",1790 => X"00000000",1791 => X"00000000",
1792 => X"00000000",1793 => X"8C510000",1794 => X"3C022000",1795 => X"34420040",
1796 => X"AC400000",1797 => X"3C032000",1798 => X"3463004C",1799 => X"3C020000",
1800 => X"24420800",1801 => X"AC620000",1802 => X"3C032000",1803 => X"34630050",
1804 => X"240200FF",1805 => X"AC620000",1806 => X"0C00001A",1807 => X"24040001",
1808 => X"3C040000",1809 => X"24841F0C",1810 => X"26310001",1811 => X"0C000080",
1812 => X"AE110000",1813 => X"02202025",1814 => X"27A50010",1815 => X"0C00019B",
1816 => X"2406000A",1817 => X"0C00008E",1818 => X"27A40010",1819 => X"0C0000C4",
1820 => X"00000000",1821 => X"00408825",1822 => X"0C0000D6",1823 => X"322400FF",
1824 => X"1000FFFA",1825 => X"00000000",1826 => X"27BDFFD0",1827 => X"AFBF0028",
1828 => X"AFB10024",1829 => X"AFB00020",1830 => X"00808825",1831 => X"0C000331",
1832 => X"27A50010",1833 => X"3C040000",1834 => X"24841EC4",1835 => X"0C000099",
1836 => X"24050003",1837 => X"8FA40010",1838 => X"3C100000",1839 => X"26101F60",
1840 => X"2402003B",1841 => X"A202000B",1842 => X"0C000261",1843 => X"02002825",
1844 => X"02002025",1845 => X"0C000099",1846 => X"2405000C",1847 => X"8FA40014",
1848 => X"0C000261",1849 => X"02002825",1850 => X"02002025",1851 => X"0C000099",
1852 => X"2405000C",1853 => X"27A40018",1854 => X"02002825",1855 => X"0C0001E7",
1856 => X"24060001",1857 => X"02002025",1858 => X"0C000099",1859 => X"24050002",
1860 => X"0C0000D6",1861 => X"2404003B",1862 => X"27A40010",1863 => X"3C050000",
1864 => X"0C000343",1865 => X"24A51F1C",1866 => X"10400019",1867 => X"24020011",
1868 => X"93A30018",1869 => X"00000000",1870 => X"14620006",1871 => X"24020001",
1872 => X"02202025",1873 => X"0C00041A",1874 => X"27A50010",1875 => X"10000010",
1876 => X"00000000",1877 => X"14620006",1878 => X"24020006",1879 => X"02202025",
1880 => X"0C0003D8",1881 => X"27A50010",1882 => X"10000009",1883 => X"00000000",
1884 => X"14620005",1885 => X"02202025",1886 => X"0C000405",1887 => X"27A50010",
1888 => X"10000003",1889 => X"00000000",1890 => X"0C000446",1891 => X"27A50010",
1892 => X"8FBF0028",1893 => X"8FB10024",1894 => X"8FB00020",1895 => X"03E00008",
1896 => X"27BD0030",1897 => X"27BDFFE8",1898 => X"AFBF0010",1899 => X"3C022001",
1900 => X"34425030",1901 => X"00A21026",1902 => X"8C420000",1903 => X"00000000",
1904 => X"3043FFFF",1905 => X"24020800",1906 => X"1062000B",1907 => X"00603025",
1908 => X"24020806",1909 => X"1062000F",1910 => X"2CC20600",1911 => X"1040000F",
1912 => X"3C02F000",1913 => X"8C860000",1914 => X"3C034000",1915 => X"00C21024",
1916 => X"14430005",1917 => X"3C020001",1918 => X"0C000722",1919 => X"00000000",
1920 => X"10000006",1921 => X"00000000",1922 => X"34420800",1923 => X"14C20003",
1924 => X"00000000",1925 => X"0C00045D",1926 => X"00000000",1927 => X"8FBF0010",
1928 => X"00000000",1929 => X"03E00008",1930 => X"27BD0018",1931 => X"00000000",
1932 => X"00000000",1933 => X"00000000",1934 => X"00000000",1935 => X"00000000",
1936 => X"00000000",1937 => X"0A0D0000",1938 => X"5A595857",1939 => X"56555453",
1940 => X"5251504F",1941 => X"4E4D4C4B",1942 => X"4A494847",1943 => X"46454443",
1944 => X"42413938",1945 => X"37363534",1946 => X"33323130",1947 => X"31323334",
1948 => X"35363738",1949 => X"39414243",1950 => X"44454647",1951 => X"48494A4B",
1952 => X"4C4D4E4F",1953 => X"50515253",1954 => X"54555657",1955 => X"58595A00",
1956 => X"30313233",1957 => X"34353637",1958 => X"38394142",1959 => X"43444546",
1960 => X"00000000",1961 => X"0A537461",1962 => X"636B6564",1963 => X"210A0000",
1964 => X"443A0000",1965 => X"433A0000",1966 => X"553A0000",1967 => X"493A0000",
1968 => X"0A410000",1969 => X"0A493A00",1970 => X"61000000",1971 => X"63000000",
1972 => X"0A495020",1973 => X"41646472",1974 => X"6573733A",1975 => X"20000000",
1976 => X"3B000000",1977 => X"4C656173",1978 => X"653A2000",1979 => X"3139322E",
1980 => X"3136382E",1981 => X"3130342E",1982 => X"36340000",1983 => X"48656C6C",
1984 => X"6F20576F",1985 => X"726C640A",1986 => X"00000000",1987 => X"48656C6C",
1988 => X"6F20576F",1989 => X"726C6420",1990 => X"00000000",1991 => X"00000001",
1992 => X"00000001",1993 => X"01000000",1994 => X"2ABCDEF0",1995 => X"20000040",
1996 => X"20000044",1997 => X"2000004C",1998 => X"20000050",1999 => X"00000000",
2000 => X"00000000",2001 => X"00000000",2002 => X"00000000",2003 => X"00000000",
2004 => X"FFFFFFFF",2005 => X"00000000",
    others => (others => '0')
    );
  signal addr_i : std_logic_vector(M-1 downto 0);

  signal din_i : std_logic_vector(N*8-1 downto 0);

  
begin  -- logic

  din_i <= to_X01(din);


  PROCESS_A : process (clk)
  begin  -- process WRITE_PROCESS
    if rising_edge(clk) then           -- rising clock edge
      addr_i <= addr;
      for i in 0 to N-1 loop
        if wbe(i) = '1' then
          ram(to_integer(unsigned(addr)))(8*i+7 downto 8*i) <= din_i(8*i+7 downto 8*i);
        end if;
      end loop;  -- i
    end if;
  end process PROCESS_A;

  dout <= ram(to_integer(unsigned(addr_i)));

end logic;
